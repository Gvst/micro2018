
module full_control_system ( clk_sm, SM1_voltage, SM1_issued_this_cycle, 
        SM1_remaining, SM2_voltage, SM2_issued_this_cycle, SM2_remaining, 
        SM3_voltage, SM3_issued_this_cycle, SM3_remaining, SM4_voltage, 
        SM4_issued_this_cycle, SM4_remaining, SM5_voltage, 
        SM5_issued_this_cycle, SM5_remaining, SM6_voltage, 
        SM6_issued_this_cycle, SM6_remaining, SM7_voltage, 
        SM7_issued_this_cycle, SM7_remaining, SM8_voltage, 
        SM8_issued_this_cycle, SM8_remaining, SM9_voltage, 
        SM9_issued_this_cycle, SM9_remaining, SM10_voltage, 
        SM10_issued_this_cycle, SM10_remaining, SM11_voltage, 
        SM11_issued_this_cycle, SM11_remaining, SM12_voltage, 
        SM12_issued_this_cycle, SM12_remaining, SM13_voltage, 
        SM13_issued_this_cycle, SM13_remaining, SM14_voltage, 
        SM14_issued_this_cycle, SM14_remaining, SM15_voltage, 
        SM15_issued_this_cycle, SM15_remaining, SM16_voltage, 
        SM16_issued_this_cycle, SM16_remaining );
  input [7:0] SM1_voltage;
  input [4:0] SM1_issued_this_cycle;
  output [4:0] SM1_remaining;
  input [7:0] SM2_voltage;
  input [4:0] SM2_issued_this_cycle;
  output [4:0] SM2_remaining;
  input [7:0] SM3_voltage;
  input [4:0] SM3_issued_this_cycle;
  output [4:0] SM3_remaining;
  input [7:0] SM4_voltage;
  input [4:0] SM4_issued_this_cycle;
  output [4:0] SM4_remaining;
  input [7:0] SM5_voltage;
  input [4:0] SM5_issued_this_cycle;
  output [4:0] SM5_remaining;
  input [7:0] SM6_voltage;
  input [4:0] SM6_issued_this_cycle;
  output [4:0] SM6_remaining;
  input [7:0] SM7_voltage;
  input [4:0] SM7_issued_this_cycle;
  output [4:0] SM7_remaining;
  input [7:0] SM8_voltage;
  input [4:0] SM8_issued_this_cycle;
  output [4:0] SM8_remaining;
  input [7:0] SM9_voltage;
  input [4:0] SM9_issued_this_cycle;
  output [4:0] SM9_remaining;
  input [7:0] SM10_voltage;
  input [4:0] SM10_issued_this_cycle;
  output [4:0] SM10_remaining;
  input [7:0] SM11_voltage;
  input [4:0] SM11_issued_this_cycle;
  output [4:0] SM11_remaining;
  input [7:0] SM12_voltage;
  input [4:0] SM12_issued_this_cycle;
  output [4:0] SM12_remaining;
  input [7:0] SM13_voltage;
  input [4:0] SM13_issued_this_cycle;
  output [4:0] SM13_remaining;
  input [7:0] SM14_voltage;
  input [4:0] SM14_issued_this_cycle;
  output [4:0] SM14_remaining;
  input [7:0] SM15_voltage;
  input [4:0] SM15_issued_this_cycle;
  output [4:0] SM15_remaining;
  input [7:0] SM16_voltage;
  input [4:0] SM16_issued_this_cycle;
  output [4:0] SM16_remaining;
  input clk_sm;
  wire   n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         clk_controller, N3, N5, N6, N11, N13, \DUT_controller/N159 ,
         \DUT_controller/N158 , \DUT_controller/N157 , \DUT_controller/N156 ,
         \DUT_controller/N155 , \DUT_controller/N149 , \DUT_controller/N148 ,
         \DUT_controller/N147 , \DUT_controller/N146 , \DUT_controller/N145 ,
         \DUT_controller/N139 , \DUT_controller/N138 , \DUT_controller/N137 ,
         \DUT_controller/N136 , \DUT_controller/N135 , \DUT_controller/N129 ,
         \DUT_controller/N128 , \DUT_controller/N127 , \DUT_controller/N126 ,
         \DUT_controller/N125 , \DUT_controller/N119 , \DUT_controller/N118 ,
         \DUT_controller/N117 , \DUT_controller/N116 , \DUT_controller/N115 ,
         \DUT_controller/N109 , \DUT_controller/N108 , \DUT_controller/N107 ,
         \DUT_controller/N106 , \DUT_controller/N105 , \DUT_controller/N99 ,
         \DUT_controller/N98 , \DUT_controller/N97 , \DUT_controller/N96 ,
         \DUT_controller/N95 , \DUT_controller/N89 , \DUT_controller/N88 ,
         \DUT_controller/N87 , \DUT_controller/N86 , \DUT_controller/N85 ,
         \DUT_controller/N79 , \DUT_controller/N78 , \DUT_controller/N77 ,
         \DUT_controller/N76 , \DUT_controller/N75 , \DUT_controller/N69 ,
         \DUT_controller/N68 , \DUT_controller/N67 , \DUT_controller/N66 ,
         \DUT_controller/N65 , \DUT_controller/N59 , \DUT_controller/N58 ,
         \DUT_controller/N57 , \DUT_controller/N56 , \DUT_controller/N55 ,
         \DUT_controller/N49 , \DUT_controller/N48 , \DUT_controller/N47 ,
         \DUT_controller/N46 , \DUT_controller/N45 , \DUT_controller/N39 ,
         \DUT_controller/N38 , \DUT_controller/N37 , \DUT_controller/N36 ,
         \DUT_controller/N35 , \DUT_controller/N29 , \DUT_controller/N28 ,
         \DUT_controller/N27 , \DUT_controller/N26 , \DUT_controller/N25 ,
         \DUT_controller/N19 , \DUT_controller/N18 , \DUT_controller/N17 ,
         \DUT_controller/N16 , \DUT_controller/N15 , \DUT_controller/N9 ,
         \DUT_controller/N8 , \DUT_controller/N7 , \DUT_controller/N6 ,
         \DUT_controller/N5 , \DUT_SM1_adjuster/N20 , \DUT_SM1_adjuster/N19 ,
         \DUT_SM1_adjuster/N18 , \DUT_SM1_adjuster/N16 ,
         \DUT_SM1_adjuster/N15 , \DUT_SM1_adjuster/N14 ,
         \DUT_SM1_adjuster/N13 , \DUT_SM1_adjuster/N12 ,
         \DUT_SM2_adjuster/N20 , \DUT_SM2_adjuster/N19 ,
         \DUT_SM2_adjuster/N18 , \DUT_SM2_adjuster/N16 ,
         \DUT_SM2_adjuster/N15 , \DUT_SM2_adjuster/N14 ,
         \DUT_SM2_adjuster/N13 , \DUT_SM2_adjuster/N12 ,
         \DUT_SM3_adjuster/N20 , \DUT_SM3_adjuster/N19 ,
         \DUT_SM3_adjuster/N18 , \DUT_SM3_adjuster/N16 ,
         \DUT_SM3_adjuster/N15 , \DUT_SM3_adjuster/N14 ,
         \DUT_SM3_adjuster/N13 , \DUT_SM3_adjuster/N12 ,
         \DUT_SM4_adjuster/N20 , \DUT_SM4_adjuster/N19 ,
         \DUT_SM4_adjuster/N18 , \DUT_SM4_adjuster/N16 ,
         \DUT_SM4_adjuster/N15 , \DUT_SM4_adjuster/N14 ,
         \DUT_SM4_adjuster/N13 , \DUT_SM4_adjuster/N12 ,
         \DUT_SM5_adjuster/N20 , \DUT_SM5_adjuster/N19 ,
         \DUT_SM5_adjuster/N18 , \DUT_SM5_adjuster/N16 ,
         \DUT_SM5_adjuster/N15 , \DUT_SM5_adjuster/N14 ,
         \DUT_SM5_adjuster/N13 , \DUT_SM5_adjuster/N12 ,
         \DUT_SM6_adjuster/N20 , \DUT_SM6_adjuster/N19 ,
         \DUT_SM6_adjuster/N18 , \DUT_SM6_adjuster/N16 ,
         \DUT_SM6_adjuster/N15 , \DUT_SM6_adjuster/N14 ,
         \DUT_SM6_adjuster/N13 , \DUT_SM6_adjuster/N12 ,
         \DUT_SM7_adjuster/N20 , \DUT_SM7_adjuster/N19 ,
         \DUT_SM7_adjuster/N18 , \DUT_SM7_adjuster/N16 ,
         \DUT_SM7_adjuster/N15 , \DUT_SM7_adjuster/N14 ,
         \DUT_SM7_adjuster/N13 , \DUT_SM7_adjuster/N12 ,
         \DUT_SM8_adjuster/N20 , \DUT_SM8_adjuster/N19 ,
         \DUT_SM8_adjuster/N18 , \DUT_SM8_adjuster/N16 ,
         \DUT_SM8_adjuster/N15 , \DUT_SM8_adjuster/N14 ,
         \DUT_SM8_adjuster/N13 , \DUT_SM8_adjuster/N12 ,
         \DUT_SM9_adjuster/N20 , \DUT_SM9_adjuster/N19 ,
         \DUT_SM9_adjuster/N18 , \DUT_SM9_adjuster/N16 ,
         \DUT_SM9_adjuster/N15 , \DUT_SM9_adjuster/N14 ,
         \DUT_SM9_adjuster/N13 , \DUT_SM9_adjuster/N12 ,
         \DUT_SM10_adjuster/N20 , \DUT_SM10_adjuster/N19 ,
         \DUT_SM10_adjuster/N18 , \DUT_SM10_adjuster/N16 ,
         \DUT_SM10_adjuster/N15 , \DUT_SM10_adjuster/N14 ,
         \DUT_SM10_adjuster/N13 , \DUT_SM10_adjuster/N12 ,
         \DUT_SM11_adjuster/N20 , \DUT_SM11_adjuster/N19 ,
         \DUT_SM11_adjuster/N18 , \DUT_SM11_adjuster/N16 ,
         \DUT_SM11_adjuster/N15 , \DUT_SM11_adjuster/N14 ,
         \DUT_SM11_adjuster/N13 , \DUT_SM11_adjuster/N12 ,
         \DUT_SM12_adjuster/N20 , \DUT_SM12_adjuster/N19 ,
         \DUT_SM12_adjuster/N18 , \DUT_SM12_adjuster/N16 ,
         \DUT_SM12_adjuster/N15 , \DUT_SM12_adjuster/N14 ,
         \DUT_SM12_adjuster/N13 , \DUT_SM12_adjuster/N12 ,
         \DUT_SM13_adjuster/N20 , \DUT_SM13_adjuster/N19 ,
         \DUT_SM13_adjuster/N18 , \DUT_SM13_adjuster/N16 ,
         \DUT_SM13_adjuster/N15 , \DUT_SM13_adjuster/N14 ,
         \DUT_SM13_adjuster/N13 , \DUT_SM13_adjuster/N12 ,
         \DUT_SM14_adjuster/N20 , \DUT_SM14_adjuster/N19 ,
         \DUT_SM14_adjuster/N18 , \DUT_SM14_adjuster/N16 ,
         \DUT_SM14_adjuster/N15 , \DUT_SM14_adjuster/N14 ,
         \DUT_SM14_adjuster/N13 , \DUT_SM14_adjuster/N12 ,
         \DUT_SM15_adjuster/N20 , \DUT_SM15_adjuster/N19 ,
         \DUT_SM15_adjuster/N18 , \DUT_SM15_adjuster/N16 ,
         \DUT_SM15_adjuster/N15 , \DUT_SM15_adjuster/N14 ,
         \DUT_SM15_adjuster/N13 , \DUT_SM15_adjuster/N12 ,
         \DUT_SM16_adjuster/N20 , \DUT_SM16_adjuster/N19 ,
         \DUT_SM16_adjuster/N18 , \DUT_SM16_adjuster/N16 ,
         \DUT_SM16_adjuster/N15 , \DUT_SM16_adjuster/N14 ,
         \DUT_SM16_adjuster/N13 , \DUT_SM16_adjuster/N12 , n195, n202, n204,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1240, n1242, n1243, n1299,
         n1308, n1310, n1311, n1315, n1316, n1317;
  wire   [4:0] SM1_issue_width_10_cycle;
  wire   [4:0] SM2_issue_width_10_cycle;
  wire   [4:0] SM3_issue_width_10_cycle;
  wire   [4:0] SM4_issue_width_10_cycle;
  wire   [4:0] SM5_issue_width_10_cycle;
  wire   [4:0] SM6_issue_width_10_cycle;
  wire   [4:0] SM7_issue_width_10_cycle;
  wire   [4:0] SM8_issue_width_10_cycle;
  wire   [4:0] SM9_issue_width_10_cycle;
  wire   [4:0] SM10_issue_width_10_cycle;
  wire   [4:0] SM11_issue_width_10_cycle;
  wire   [4:0] SM12_issue_width_10_cycle;
  wire   [4:0] SM13_issue_width_10_cycle;
  wire   [4:0] SM14_issue_width_10_cycle;
  wire   [4:0] SM15_issue_width_10_cycle;
  wire   [4:0] SM16_issue_width_10_cycle;
  wire   [5:0] counter;
  wire   [3:0] \DUT_SM1_adjuster/rst ;
  wire   [3:0] \DUT_SM2_adjuster/rst ;
  wire   [3:0] \DUT_SM3_adjuster/rst ;
  wire   [3:0] \DUT_SM4_adjuster/rst ;
  wire   [3:0] \DUT_SM5_adjuster/rst ;
  wire   [3:0] \DUT_SM6_adjuster/rst ;
  wire   [3:0] \DUT_SM7_adjuster/rst ;
  wire   [3:0] \DUT_SM8_adjuster/rst ;
  wire   [3:0] \DUT_SM9_adjuster/rst ;
  wire   [3:0] \DUT_SM10_adjuster/rst ;
  wire   [3:0] \DUT_SM11_adjuster/rst ;
  wire   [3:0] \DUT_SM12_adjuster/rst ;
  wire   [3:0] \DUT_SM13_adjuster/rst ;
  wire   [3:0] \DUT_SM14_adjuster/rst ;
  wire   [3:0] \DUT_SM15_adjuster/rst ;
  wire   [3:0] \DUT_SM16_adjuster/rst ;

  DFFQ_X1M_A9TR clk_controller_reg ( .D(n195), .CK(clk_sm), .Q(clk_controller)
         );
  DFFQ_X1M_A9TR \DUT_SM16_adjuster/rst_reg[0]  ( .D(n1315), .CK(clk_sm), .Q(
        \DUT_SM16_adjuster/rst [0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM8_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N76 ), .CK(clk_controller), .Q(
        SM8_issue_width_10_cycle[1]) );
  DFFQ_X1M_A9TR \DUT_controller/SM8_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N77 ), .CK(clk_controller), .Q(
        SM8_issue_width_10_cycle[2]) );
  DFFQ_X1M_A9TR \DUT_controller/SM8_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N78 ), .CK(clk_controller), .Q(
        SM8_issue_width_10_cycle[3]) );
  DFFQ_X1M_A9TR \DUT_controller/SM8_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N79 ), .CK(clk_controller), .Q(
        SM8_issue_width_10_cycle[4]) );
  DFFQ_X1M_A9TR \DUT_controller/SM7_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N66 ), .CK(clk_controller), .Q(
        SM7_issue_width_10_cycle[1]) );
  DFFQ_X1M_A9TR \DUT_controller/SM7_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N67 ), .CK(clk_controller), .Q(
        SM7_issue_width_10_cycle[2]) );
  DFFQ_X1M_A9TR \DUT_controller/SM7_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N68 ), .CK(clk_controller), .Q(
        SM7_issue_width_10_cycle[3]) );
  DFFQ_X1M_A9TR \DUT_controller/SM16_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N156 ), .CK(n1317), .Q(SM16_issue_width_10_cycle[1])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM16_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N157 ), .CK(n1317), .Q(SM16_issue_width_10_cycle[2])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM16_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N158 ), .CK(n1317), .Q(SM16_issue_width_10_cycle[3])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM16_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N159 ), .CK(n1317), .Q(SM16_issue_width_10_cycle[4])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM15_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N146 ), .CK(n1317), .Q(SM15_issue_width_10_cycle[1])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM15_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N147 ), .CK(n1317), .Q(SM15_issue_width_10_cycle[2])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM15_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N148 ), .CK(n1317), .Q(SM15_issue_width_10_cycle[3])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM15_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N149 ), .CK(n1317), .Q(SM15_issue_width_10_cycle[4])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM14_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N136 ), .CK(n1317), .Q(SM14_issue_width_10_cycle[1])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM14_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N137 ), .CK(n1317), .Q(SM14_issue_width_10_cycle[2])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM14_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N138 ), .CK(n1317), .Q(SM14_issue_width_10_cycle[3])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM14_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N139 ), .CK(n1317), .Q(SM14_issue_width_10_cycle[4])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM13_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N126 ), .CK(n1317), .Q(SM13_issue_width_10_cycle[1])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM13_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N127 ), .CK(n1317), .Q(SM13_issue_width_10_cycle[2])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM13_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N128 ), .CK(n1317), .Q(SM13_issue_width_10_cycle[3])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM13_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N129 ), .CK(n1317), .Q(SM13_issue_width_10_cycle[4])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM3_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N27 ), .CK(n1317), .Q(SM3_issue_width_10_cycle[2]) );
  DFFQ_X1M_A9TR \DUT_controller/SM3_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N29 ), .CK(n1317), .Q(SM3_issue_width_10_cycle[4]) );
  DFFQ_X1M_A9TR \DUT_controller/SM2_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N16 ), .CK(n1317), .Q(SM2_issue_width_10_cycle[1]) );
  DFFQ_X1M_A9TR \DUT_controller/SM2_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N18 ), .CK(n1317), .Q(SM2_issue_width_10_cycle[3]) );
  DFFQ_X1M_A9TR \DUT_controller/SM12_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N116 ), .CK(n1317), .Q(SM12_issue_width_10_cycle[1])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM12_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N117 ), .CK(n1317), .Q(SM12_issue_width_10_cycle[2])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM12_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N118 ), .CK(n1317), .Q(SM12_issue_width_10_cycle[3])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM12_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N119 ), .CK(n1317), .Q(SM12_issue_width_10_cycle[4])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM11_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N106 ), .CK(n1317), .Q(SM11_issue_width_10_cycle[1])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM11_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N107 ), .CK(n1317), .Q(SM11_issue_width_10_cycle[2])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM11_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N108 ), .CK(n1317), .Q(SM11_issue_width_10_cycle[3])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM11_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N109 ), .CK(n1317), .Q(SM11_issue_width_10_cycle[4])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM10_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N96 ), .CK(n1317), .Q(SM10_issue_width_10_cycle[1]) );
  DFFQ_X1M_A9TR \DUT_controller/SM10_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N97 ), .CK(n1317), .Q(SM10_issue_width_10_cycle[2]) );
  DFFQ_X1M_A9TR \DUT_controller/SM10_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N98 ), .CK(n1317), .Q(SM10_issue_width_10_cycle[3]) );
  DFFQ_X1M_A9TR \DUT_controller/SM10_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N99 ), .CK(n1317), .Q(SM10_issue_width_10_cycle[4]) );
  DFFQ_X1M_A9TR \DUT_controller/SM9_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N86 ), .CK(n1317), .Q(SM9_issue_width_10_cycle[1]) );
  DFFQ_X1M_A9TR \DUT_controller/SM9_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N87 ), .CK(n1317), .Q(SM9_issue_width_10_cycle[2]) );
  DFFQ_X1M_A9TR \DUT_controller/SM9_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N88 ), .CK(n1317), .Q(SM9_issue_width_10_cycle[3]) );
  DFFQ_X1M_A9TR \DUT_controller/SM9_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N89 ), .CK(n1317), .Q(SM9_issue_width_10_cycle[4]) );
  DFFQ_X1M_A9TR \DUT_controller/SM7_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N69 ), .CK(n1317), .Q(SM7_issue_width_10_cycle[4]) );
  DFFQ_X1M_A9TR \DUT_controller/SM6_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N56 ), .CK(n1317), .Q(SM6_issue_width_10_cycle[1]) );
  DFFQ_X1M_A9TR \DUT_controller/SM6_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N57 ), .CK(n1317), .Q(SM6_issue_width_10_cycle[2]) );
  DFFQ_X1M_A9TR \DUT_controller/SM6_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N58 ), .CK(n1317), .Q(SM6_issue_width_10_cycle[3]) );
  DFFQ_X1M_A9TR \DUT_controller/SM6_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N59 ), .CK(n1317), .Q(SM6_issue_width_10_cycle[4]) );
  DFFQ_X1M_A9TR \DUT_controller/SM5_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N46 ), .CK(n1317), .Q(SM5_issue_width_10_cycle[1]) );
  DFFQ_X1M_A9TR \DUT_controller/SM5_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N47 ), .CK(n1317), .Q(SM5_issue_width_10_cycle[2]) );
  DFFQ_X1M_A9TR \DUT_controller/SM5_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N48 ), .CK(n1317), .Q(SM5_issue_width_10_cycle[3]) );
  DFFQ_X1M_A9TR \DUT_controller/SM5_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N49 ), .CK(n1317), .Q(SM5_issue_width_10_cycle[4]) );
  DFFQ_X1M_A9TR \DUT_controller/SM4_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N36 ), .CK(n1317), .Q(SM4_issue_width_10_cycle[1]) );
  DFFQ_X1M_A9TR \DUT_controller/SM4_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N37 ), .CK(n1317), .Q(SM4_issue_width_10_cycle[2]) );
  DFFQ_X1M_A9TR \DUT_controller/SM4_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N38 ), .CK(n1317), .Q(SM4_issue_width_10_cycle[3]) );
  DFFQ_X1M_A9TR \DUT_controller/SM4_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N39 ), .CK(n1317), .Q(SM4_issue_width_10_cycle[4]) );
  DFFQ_X1M_A9TR \DUT_controller/SM3_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N26 ), .CK(n1317), .Q(SM3_issue_width_10_cycle[1]) );
  DFFQ_X1M_A9TR \DUT_controller/SM3_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N28 ), .CK(n1317), .Q(SM3_issue_width_10_cycle[3]) );
  DFFQ_X1M_A9TR \DUT_controller/SM2_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N17 ), .CK(n1317), .Q(SM2_issue_width_10_cycle[2]) );
  DFFQ_X1M_A9TR \DUT_controller/SM2_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N19 ), .CK(n1317), .Q(SM2_issue_width_10_cycle[4]) );
  DFFQ_X1M_A9TR \DUT_controller/SM1_issue_width_10_cycle_reg[1]  ( .D(
        \DUT_controller/N6 ), .CK(n1317), .Q(SM1_issue_width_10_cycle[1]) );
  DFFQ_X1M_A9TR \DUT_controller/SM1_issue_width_10_cycle_reg[2]  ( .D(
        \DUT_controller/N7 ), .CK(n1317), .Q(SM1_issue_width_10_cycle[2]) );
  DFFQ_X1M_A9TR \DUT_controller/SM1_issue_width_10_cycle_reg[3]  ( .D(
        \DUT_controller/N8 ), .CK(n1317), .Q(SM1_issue_width_10_cycle[3]) );
  DFFQ_X1M_A9TR \DUT_controller/SM1_issue_width_10_cycle_reg[4]  ( .D(
        \DUT_controller/N9 ), .CK(n1317), .Q(SM1_issue_width_10_cycle[4]) );
  DFFQ_X1M_A9TR \DUT_controller/SM16_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N155 ), .CK(clk_controller), .Q(
        SM16_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM7_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N65 ), .CK(clk_controller), .Q(
        SM7_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM15_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N145 ), .CK(n1317), .Q(SM15_issue_width_10_cycle[0])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM14_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N135 ), .CK(n1317), .Q(SM14_issue_width_10_cycle[0])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM13_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N125 ), .CK(n1317), .Q(SM13_issue_width_10_cycle[0])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM12_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N115 ), .CK(n1317), .Q(SM12_issue_width_10_cycle[0])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM3_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N25 ), .CK(n1317), .Q(SM3_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM1_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N5 ), .CK(n1317), .Q(SM1_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM11_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N105 ), .CK(n1317), .Q(SM11_issue_width_10_cycle[0])
         );
  DFFQ_X1M_A9TR \DUT_controller/SM10_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N95 ), .CK(n1317), .Q(SM10_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM9_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N85 ), .CK(n1317), .Q(SM9_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM8_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N75 ), .CK(n1317), .Q(SM8_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM6_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N55 ), .CK(n1317), .Q(SM6_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM5_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N45 ), .CK(n1317), .Q(SM5_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM4_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N35 ), .CK(n1317), .Q(SM4_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \DUT_controller/SM2_issue_width_10_cycle_reg[0]  ( .D(
        \DUT_controller/N15 ), .CK(n1317), .Q(SM2_issue_width_10_cycle[0]) );
  DFFQ_X1M_A9TR \counter_reg[5]  ( .D(N6), .CK(clk_sm), .Q(counter[5]) );
  DFFQ_X1M_A9TR \counter_reg[4]  ( .D(N5), .CK(clk_sm), .Q(counter[4]) );
  DFFQ_X1M_A9TR \counter_reg[3]  ( .D(N13), .CK(clk_sm), .Q(counter[3]) );
  DFFQ_X1M_A9TR \counter_reg[2]  ( .D(N3), .CK(clk_sm), .Q(counter[2]) );
  DFFQ_X1M_A9TR \counter_reg[1]  ( .D(N11), .CK(clk_sm), .Q(counter[1]) );
  DFFQ_X1M_A9TR \DUT_SM1_adjuster/rst_reg[2]  ( .D(\DUT_SM1_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM1_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM2_adjuster/rst_reg[2]  ( .D(\DUT_SM2_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM2_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM3_adjuster/rst_reg[2]  ( .D(\DUT_SM3_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM3_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM4_adjuster/rst_reg[2]  ( .D(\DUT_SM4_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM4_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM5_adjuster/rst_reg[2]  ( .D(\DUT_SM5_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM5_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM6_adjuster/rst_reg[2]  ( .D(\DUT_SM6_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM6_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM7_adjuster/rst_reg[2]  ( .D(\DUT_SM7_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM7_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM8_adjuster/rst_reg[2]  ( .D(\DUT_SM8_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM8_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM9_adjuster/rst_reg[2]  ( .D(\DUT_SM9_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM9_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM10_adjuster/rst_reg[2]  ( .D(\DUT_SM10_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM10_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM11_adjuster/rst_reg[2]  ( .D(\DUT_SM11_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM11_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM12_adjuster/rst_reg[2]  ( .D(\DUT_SM12_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM12_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM13_adjuster/rst_reg[2]  ( .D(\DUT_SM13_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM13_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM14_adjuster/rst_reg[2]  ( .D(\DUT_SM14_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM14_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM15_adjuster/rst_reg[2]  ( .D(\DUT_SM15_adjuster/N19 ), 
        .CK(clk_sm), .Q(\DUT_SM15_adjuster/rst [2]) );
  DFFQ_X1M_A9TR \DUT_SM1_adjuster/rst_reg[1]  ( .D(\DUT_SM1_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM1_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM2_adjuster/rst_reg[1]  ( .D(\DUT_SM2_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM2_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM3_adjuster/rst_reg[1]  ( .D(\DUT_SM3_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM3_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM4_adjuster/rst_reg[1]  ( .D(\DUT_SM4_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM4_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM5_adjuster/rst_reg[1]  ( .D(\DUT_SM5_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM5_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM6_adjuster/rst_reg[1]  ( .D(\DUT_SM6_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM6_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM7_adjuster/rst_reg[1]  ( .D(\DUT_SM7_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM7_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM8_adjuster/rst_reg[1]  ( .D(\DUT_SM8_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM8_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM9_adjuster/rst_reg[1]  ( .D(\DUT_SM9_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM9_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM10_adjuster/rst_reg[1]  ( .D(\DUT_SM10_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM10_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM11_adjuster/rst_reg[1]  ( .D(\DUT_SM11_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM11_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM12_adjuster/rst_reg[1]  ( .D(\DUT_SM12_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM12_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM13_adjuster/rst_reg[1]  ( .D(\DUT_SM13_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM13_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM14_adjuster/rst_reg[1]  ( .D(\DUT_SM14_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM14_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM15_adjuster/rst_reg[1]  ( .D(\DUT_SM15_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM15_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM16_adjuster/rst_reg[1]  ( .D(\DUT_SM16_adjuster/N18 ), 
        .CK(clk_sm), .Q(\DUT_SM16_adjuster/rst [1]) );
  DFFQ_X1M_A9TR \DUT_SM1_adjuster/rst_reg[3]  ( .D(\DUT_SM1_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM1_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM2_adjuster/rst_reg[3]  ( .D(\DUT_SM2_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM2_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM3_adjuster/rst_reg[3]  ( .D(\DUT_SM3_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM3_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM4_adjuster/rst_reg[3]  ( .D(\DUT_SM4_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM4_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM5_adjuster/rst_reg[3]  ( .D(\DUT_SM5_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM5_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM6_adjuster/rst_reg[3]  ( .D(\DUT_SM6_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM6_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM7_adjuster/rst_reg[3]  ( .D(\DUT_SM7_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM7_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM8_adjuster/rst_reg[3]  ( .D(\DUT_SM8_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM8_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM9_adjuster/rst_reg[3]  ( .D(\DUT_SM9_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM9_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM10_adjuster/rst_reg[3]  ( .D(\DUT_SM10_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM10_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM11_adjuster/rst_reg[3]  ( .D(\DUT_SM11_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM11_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM12_adjuster/rst_reg[3]  ( .D(\DUT_SM12_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM12_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM13_adjuster/rst_reg[3]  ( .D(\DUT_SM13_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM13_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM14_adjuster/rst_reg[3]  ( .D(\DUT_SM14_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM14_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM15_adjuster/rst_reg[3]  ( .D(\DUT_SM15_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM15_adjuster/rst [3]) );
  DFFQ_X1M_A9TR \DUT_SM16_adjuster/rst_reg[3]  ( .D(\DUT_SM16_adjuster/N20 ), 
        .CK(clk_sm), .Q(\DUT_SM16_adjuster/rst [3]) );
  DFFQN_X1M_A9TR \DUT_SM16_adjuster/rst_reg[2]  ( .D(\DUT_SM16_adjuster/N19 ), 
        .CK(clk_sm), .QN(n1316) );
  DFFQ_X4M_A9TR \DUT_SM16_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM16_adjuster/N14 ), .CK(clk_sm), .Q(n1395) );
  DFFQ_X4M_A9TR \DUT_SM15_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM15_adjuster/N14 ), .CK(clk_sm), .Q(n1390) );
  DFFQ_X4M_A9TR \DUT_SM14_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM14_adjuster/N14 ), .CK(clk_sm), .Q(n1385) );
  DFFQ_X4M_A9TR \DUT_SM13_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM13_adjuster/N14 ), .CK(clk_sm), .Q(n1380) );
  DFFQ_X4M_A9TR \DUT_SM10_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM10_adjuster/N14 ), .CK(clk_sm), .Q(n1365) );
  DFFQ_X4M_A9TR \DUT_SM9_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM9_adjuster/N14 ), .CK(clk_sm), .Q(n1360) );
  DFFQ_X4M_A9TR \DUT_SM12_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM12_adjuster/N14 ), .CK(clk_sm), .Q(n1375) );
  DFFQ_X4M_A9TR \DUT_SM11_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM11_adjuster/N14 ), .CK(clk_sm), .Q(n1370) );
  DFFQ_X4M_A9TR \DUT_SM7_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM7_adjuster/N14 ), .CK(clk_sm), .Q(n1350) );
  DFFQ_X4M_A9TR \DUT_SM6_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM6_adjuster/N14 ), .CK(clk_sm), .Q(n1345) );
  DFFQ_X4M_A9TR \DUT_SM5_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM5_adjuster/N14 ), .CK(clk_sm), .Q(n1340) );
  DFFQ_X4M_A9TR \DUT_SM2_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM2_adjuster/N14 ), .CK(clk_sm), .Q(n1325) );
  DFFQ_X4M_A9TR \DUT_SM1_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM1_adjuster/N14 ), .CK(clk_sm), .Q(n1320) );
  DFFQ_X4M_A9TR \DUT_SM8_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM8_adjuster/N14 ), .CK(clk_sm), .Q(n1355) );
  DFFQ_X4M_A9TR \DUT_SM4_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM4_adjuster/N14 ), .CK(clk_sm), .Q(n1335) );
  DFFQ_X4M_A9TR \DUT_SM3_adjuster/remaining_reg[2]  ( .D(
        \DUT_SM3_adjuster/N14 ), .CK(clk_sm), .Q(n1330) );
  DFFQ_X4M_A9TR \DUT_SM5_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM5_adjuster/N12 ), .CK(clk_sm), .Q(n1342) );
  DFFQ_X4M_A9TR \DUT_SM12_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM12_adjuster/N12 ), .CK(clk_sm), .Q(n1377) );
  DFFQ_X4M_A9TR \DUT_SM10_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM10_adjuster/N12 ), .CK(clk_sm), .Q(n1367) );
  DFFQ_X2M_A9TR \DUT_SM2_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM2_adjuster/N13 ), .CK(clk_sm), .Q(n1326) );
  DFFQ_X2M_A9TR \DUT_SM1_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM1_adjuster/N13 ), .CK(clk_sm), .Q(n1321) );
  DFFQ_X2M_A9TR \DUT_SM6_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM6_adjuster/N13 ), .CK(clk_sm), .Q(n1346) );
  DFFQ_X2M_A9TR \DUT_SM5_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM5_adjuster/N13 ), .CK(clk_sm), .Q(n1341) );
  DFFQ_X2M_A9TR \DUT_SM4_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM4_adjuster/N13 ), .CK(clk_sm), .Q(n1336) );
  DFFQ_X2M_A9TR \DUT_SM3_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM3_adjuster/N13 ), .CK(clk_sm), .Q(n1331) );
  DFFQ_X2M_A9TR \DUT_SM10_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM10_adjuster/N13 ), .CK(clk_sm), .Q(n1366) );
  DFFQ_X2M_A9TR \DUT_SM9_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM9_adjuster/N13 ), .CK(clk_sm), .Q(n1361) );
  DFFQ_X2M_A9TR \DUT_SM8_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM8_adjuster/N13 ), .CK(clk_sm), .Q(n1356) );
  DFFQ_X2M_A9TR \DUT_SM7_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM7_adjuster/N13 ), .CK(clk_sm), .Q(n1351) );
  DFFQ_X2M_A9TR \DUT_SM14_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM14_adjuster/N13 ), .CK(clk_sm), .Q(n1386) );
  DFFQ_X2M_A9TR \DUT_SM13_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM13_adjuster/N13 ), .CK(clk_sm), .Q(n1381) );
  DFFQ_X2M_A9TR \DUT_SM12_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM12_adjuster/N13 ), .CK(clk_sm), .Q(n1376) );
  DFFQ_X2M_A9TR \DUT_SM11_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM11_adjuster/N13 ), .CK(clk_sm), .Q(n1371) );
  DFFQ_X2M_A9TR \DUT_SM16_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM16_adjuster/N13 ), .CK(clk_sm), .Q(n1396) );
  DFFQ_X2M_A9TR \DUT_SM15_adjuster/remaining_reg[1]  ( .D(
        \DUT_SM15_adjuster/N13 ), .CK(clk_sm), .Q(n1391) );
  DFFQ_X3M_A9TR \DUT_SM13_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM13_adjuster/N12 ), .CK(clk_sm), .Q(n1382) );
  DFFQ_X3M_A9TR \DUT_SM9_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM9_adjuster/N12 ), .CK(clk_sm), .Q(n1362) );
  DFFQ_X3M_A9TR \DUT_SM16_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM16_adjuster/N12 ), .CK(clk_sm), .Q(n1397) );
  DFFQ_X3M_A9TR \DUT_SM15_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM15_adjuster/N12 ), .CK(clk_sm), .Q(n1392) );
  DFFQ_X3M_A9TR \DUT_SM14_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM14_adjuster/N12 ), .CK(clk_sm), .Q(n1387) );
  DFFQ_X3M_A9TR \DUT_SM11_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM11_adjuster/N12 ), .CK(clk_sm), .Q(n1372) );
  DFFQ_X3M_A9TR \DUT_SM6_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM6_adjuster/N12 ), .CK(clk_sm), .Q(n1347) );
  DFFQ_X3M_A9TR \DUT_SM2_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM2_adjuster/N12 ), .CK(clk_sm), .Q(n1327) );
  DFFQ_X3M_A9TR \DUT_SM1_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM1_adjuster/N12 ), .CK(clk_sm), .Q(n1322) );
  DFFQ_X3M_A9TR \DUT_SM8_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM8_adjuster/N12 ), .CK(clk_sm), .Q(n1357) );
  DFFQ_X3M_A9TR \DUT_SM7_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM7_adjuster/N12 ), .CK(clk_sm), .Q(n1352) );
  DFFQ_X3M_A9TR \DUT_SM4_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM4_adjuster/N12 ), .CK(clk_sm), .Q(n1337) );
  DFFQ_X3M_A9TR \DUT_SM3_adjuster/remaining_reg[0]  ( .D(
        \DUT_SM3_adjuster/N12 ), .CK(clk_sm), .Q(n1332) );
  DFFQ_X2M_A9TR \DUT_SM2_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM2_adjuster/N15 ), .CK(clk_sm), .Q(n1324) );
  DFFQ_X2M_A9TR \DUT_SM1_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM1_adjuster/N15 ), .CK(clk_sm), .Q(n1319) );
  DFFQ_X2M_A9TR \DUT_SM6_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM6_adjuster/N15 ), .CK(clk_sm), .Q(n1344) );
  DFFQ_X2M_A9TR \DUT_SM5_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM5_adjuster/N15 ), .CK(clk_sm), .Q(n1339) );
  DFFQ_X2M_A9TR \DUT_SM4_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM4_adjuster/N15 ), .CK(clk_sm), .Q(n1334) );
  DFFQ_X2M_A9TR \DUT_SM3_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM3_adjuster/N15 ), .CK(clk_sm), .Q(n1329) );
  DFFQ_X2M_A9TR \DUT_SM10_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM10_adjuster/N15 ), .CK(clk_sm), .Q(n1364) );
  DFFQ_X2M_A9TR \DUT_SM9_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM9_adjuster/N15 ), .CK(clk_sm), .Q(n1359) );
  DFFQ_X2M_A9TR \DUT_SM8_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM8_adjuster/N15 ), .CK(clk_sm), .Q(n1354) );
  DFFQ_X2M_A9TR \DUT_SM7_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM7_adjuster/N15 ), .CK(clk_sm), .Q(n1349) );
  DFFQ_X2M_A9TR \DUT_SM14_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM14_adjuster/N15 ), .CK(clk_sm), .Q(n1384) );
  DFFQ_X2M_A9TR \DUT_SM13_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM13_adjuster/N15 ), .CK(clk_sm), .Q(n1379) );
  DFFQ_X2M_A9TR \DUT_SM12_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM12_adjuster/N15 ), .CK(clk_sm), .Q(n1374) );
  DFFQ_X2M_A9TR \DUT_SM11_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM11_adjuster/N15 ), .CK(clk_sm), .Q(n1369) );
  DFFQ_X2M_A9TR \DUT_SM16_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM16_adjuster/N15 ), .CK(clk_sm), .Q(n1394) );
  DFFQ_X2M_A9TR \DUT_SM15_adjuster/remaining_reg[3]  ( .D(
        \DUT_SM15_adjuster/N15 ), .CK(clk_sm), .Q(n1389) );
  DFFQ_X2M_A9TR \DUT_SM2_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM2_adjuster/N16 ), .CK(clk_sm), .Q(n1323) );
  DFFQ_X2M_A9TR \DUT_SM1_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM1_adjuster/N16 ), .CK(clk_sm), .Q(n1318) );
  DFFQ_X2M_A9TR \DUT_SM6_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM6_adjuster/N16 ), .CK(clk_sm), .Q(n1343) );
  DFFQ_X2M_A9TR \DUT_SM5_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM5_adjuster/N16 ), .CK(clk_sm), .Q(n1338) );
  DFFQ_X2M_A9TR \DUT_SM4_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM4_adjuster/N16 ), .CK(clk_sm), .Q(n1333) );
  DFFQ_X2M_A9TR \DUT_SM3_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM3_adjuster/N16 ), .CK(clk_sm), .Q(n1328) );
  DFFQ_X2M_A9TR \DUT_SM10_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM10_adjuster/N16 ), .CK(clk_sm), .Q(n1363) );
  DFFQ_X2M_A9TR \DUT_SM9_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM9_adjuster/N16 ), .CK(clk_sm), .Q(n1358) );
  DFFQ_X2M_A9TR \DUT_SM8_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM8_adjuster/N16 ), .CK(clk_sm), .Q(n1353) );
  DFFQ_X2M_A9TR \DUT_SM7_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM7_adjuster/N16 ), .CK(clk_sm), .Q(n1348) );
  DFFQ_X2M_A9TR \DUT_SM14_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM14_adjuster/N16 ), .CK(clk_sm), .Q(n1383) );
  DFFQ_X2M_A9TR \DUT_SM13_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM13_adjuster/N16 ), .CK(clk_sm), .Q(n1378) );
  DFFQ_X2M_A9TR \DUT_SM12_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM12_adjuster/N16 ), .CK(clk_sm), .Q(n1373) );
  DFFQ_X2M_A9TR \DUT_SM11_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM11_adjuster/N16 ), .CK(clk_sm), .Q(n1368) );
  DFFQ_X2M_A9TR \DUT_SM16_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM16_adjuster/N16 ), .CK(clk_sm), .Q(n1393) );
  DFFQ_X2M_A9TR \DUT_SM15_adjuster/remaining_reg[4]  ( .D(
        \DUT_SM15_adjuster/N16 ), .CK(clk_sm), .Q(n1388) );
  BUFH_X1M_A9TR U410 ( .A(n1367), .Y(n1240) );
  BUFH_X1M_A9TR U411 ( .A(n1377), .Y(n1242) );
  BUFH_X1M_A9TR U412 ( .A(n1342), .Y(n1243) );
  BUFH_X1M_A9TR U413 ( .A(n1380), .Y(n1311) );
  BUFH_X1M_A9TR U414 ( .A(n1365), .Y(n1308) );
  BUFH_X1M_A9TR U415 ( .A(n1375), .Y(n1310) );
  BUFH_X1M_A9TR U416 ( .A(n1320), .Y(n1299) );
  BUFH_X1M_A9TR U417 ( .A(n1340), .Y(n202) );
  BUFH_X1M_A9TR U418 ( .A(n1360), .Y(n204) );
  BUFH_X1M_A9TR U419 ( .A(n1395), .Y(n207) );
  BUFH_X11M_A9TR U420 ( .A(n1367), .Y(SM10_remaining[0]) );
  BUFH_X11M_A9TR U421 ( .A(n1377), .Y(SM12_remaining[0]) );
  BUFH_X11M_A9TR U422 ( .A(n1342), .Y(SM5_remaining[0]) );
  BUFH_X11M_A9TR U423 ( .A(n1320), .Y(SM1_remaining[2]) );
  BUFH_X11M_A9TR U424 ( .A(n1375), .Y(SM12_remaining[2]) );
  BUFH_X11M_A9TR U425 ( .A(n1365), .Y(SM10_remaining[2]) );
  BUFH_X11M_A9TR U426 ( .A(n1380), .Y(SM13_remaining[2]) );
  BUFH_X1M_A9TR U427 ( .A(n1380), .Y(n795) );
  INV_X0P7M_A9TR U428 ( .A(n794), .Y(n799) );
  INV_X0P7M_A9TR U429 ( .A(n800), .Y(n804) );
  INV_X0P7M_A9TR U430 ( .A(n805), .Y(n809) );
  INV_X0P7M_A9TR U431 ( .A(n810), .Y(n814) );
  INV_X0P7M_A9TR U432 ( .A(n772), .Y(n776) );
  BUFH_X1M_A9TR U433 ( .A(n1365), .Y(n778) );
  INV_X0P7M_A9TR U434 ( .A(n777), .Y(n782) );
  INV_X0P7M_A9TR U435 ( .A(n783), .Y(n787) );
  BUFH_X1M_A9TR U436 ( .A(n1375), .Y(n789) );
  INV_X0P7M_A9TR U437 ( .A(n788), .Y(n793) );
  INV_X0P7M_A9TR U438 ( .A(n815), .Y(n819) );
  INV_X0P7M_A9TR U439 ( .A(n820), .Y(n824) );
  INV_X0P7M_A9TR U440 ( .A(n762), .Y(n766) );
  INV_X0P7M_A9TR U441 ( .A(n767), .Y(n771) );
  BUFH_X1M_A9TR U442 ( .A(n1320), .Y(n841) );
  INV_X0P7M_A9TR U443 ( .A(n840), .Y(n845) );
  INV_X0P7M_A9TR U444 ( .A(n825), .Y(n829) );
  INV_X0P7M_A9TR U445 ( .A(n830), .Y(n834) );
  INV_X0P7M_A9TR U446 ( .A(n835), .Y(n839) );
  INV_X0P7M_A9TR U447 ( .A(n1381), .Y(n847) );
  NOR2_X0P7A_A9TR U448 ( .A(n738), .B(n1382), .Y(n851) );
  INV_X0P7M_A9TR U449 ( .A(n1386), .Y(n931) );
  NOR2_X0P7A_A9TR U450 ( .A(n736), .B(n1387), .Y(n935) );
  INV_X0P7M_A9TR U451 ( .A(n1391), .Y(n925) );
  NOR2_X0P7A_A9TR U452 ( .A(n734), .B(n1392), .Y(n929) );
  INV_X0P7M_A9TR U453 ( .A(n1396), .Y(n937) );
  NOR2_X0P7A_A9TR U454 ( .A(n760), .B(n1397), .Y(n941) );
  INV_X0P7M_A9TR U455 ( .A(n1361), .Y(n871) );
  NOR2_X0P7A_A9TR U456 ( .A(n746), .B(n1362), .Y(n875) );
  INV_X0P7M_A9TR U457 ( .A(n1366), .Y(n865) );
  NOR2_X0P7A_A9TR U458 ( .A(n744), .B(n256), .Y(n869) );
  INV_X0P7M_A9TR U459 ( .A(n1371), .Y(n859) );
  NOR2_X0P7A_A9TR U460 ( .A(n742), .B(n1372), .Y(n863) );
  INV_X0P7M_A9TR U461 ( .A(n1376), .Y(n853) );
  NOR2_X0P7A_A9TR U462 ( .A(n740), .B(n267), .Y(n857) );
  INV_X0P7M_A9TR U463 ( .A(n1341), .Y(n895) );
  NOR2_X0P7A_A9TR U464 ( .A(n754), .B(n228), .Y(n899) );
  INV_X0P7M_A9TR U465 ( .A(n1346), .Y(n889) );
  NOR2_X0P7A_A9TR U466 ( .A(n752), .B(n1347), .Y(n893) );
  INV_X0P7M_A9TR U467 ( .A(n1351), .Y(n883) );
  NOR2_X0P7A_A9TR U468 ( .A(n750), .B(n1352), .Y(n887) );
  INV_X0P7M_A9TR U469 ( .A(n1356), .Y(n877) );
  NOR2_X0P7A_A9TR U470 ( .A(n748), .B(n1357), .Y(n881) );
  INV_X0P7M_A9TR U471 ( .A(n1321), .Y(n919) );
  NOR2_X0P7A_A9TR U472 ( .A(n732), .B(n1322), .Y(n923) );
  INV_X0P7M_A9TR U473 ( .A(n1326), .Y(n913) );
  NOR2_X0P7A_A9TR U474 ( .A(n730), .B(n1327), .Y(n917) );
  INV_X0P7M_A9TR U475 ( .A(n1331), .Y(n907) );
  NOR2_X0P7A_A9TR U476 ( .A(n758), .B(n1332), .Y(n911) );
  INV_X0P7M_A9TR U477 ( .A(n1336), .Y(n901) );
  NOR2_X0P7A_A9TR U478 ( .A(n756), .B(n1337), .Y(n905) );
  INV_X0P7M_A9TR U479 ( .A(n1379), .Y(n999) );
  CGENI_X1M_A9TR U480 ( .A(n1380), .B(n273), .CI(n794), .CON(n1004) );
  INV_X0P7M_A9TR U481 ( .A(n1384), .Y(n992) );
  CGENI_X1M_A9TR U482 ( .A(n1385), .B(n278), .CI(n800), .CON(n997) );
  INV_X0P7M_A9TR U483 ( .A(n1389), .Y(n985) );
  CGENI_X1M_A9TR U484 ( .A(n1390), .B(n283), .CI(n805), .CON(n990) );
  INV_X0P7M_A9TR U485 ( .A(n1394), .Y(n978) );
  CGENI_X1M_A9TR U486 ( .A(n289), .B(n288), .CI(n810), .CON(n983) );
  INV_X0P7M_A9TR U487 ( .A(n1359), .Y(n1027) );
  CGENI_X1M_A9TR U488 ( .A(n251), .B(n250), .CI(n772), .CON(n1032) );
  INV_X0P7M_A9TR U489 ( .A(n1364), .Y(n1020) );
  CGENI_X1M_A9TR U490 ( .A(n1365), .B(n257), .CI(n777), .CON(n1025) );
  INV_X0P7M_A9TR U491 ( .A(n1369), .Y(n1013) );
  CGENI_X1M_A9TR U492 ( .A(n1370), .B(n262), .CI(n783), .CON(n1018) );
  INV_X0P7M_A9TR U493 ( .A(n1374), .Y(n1006) );
  CGENI_X1M_A9TR U494 ( .A(n1375), .B(n268), .CI(n788), .CON(n1011) );
  INV_X0P7M_A9TR U495 ( .A(n1339), .Y(n971) );
  CGENI_X1M_A9TR U496 ( .A(n230), .B(n229), .CI(n815), .CON(n976) );
  INV_X0P7M_A9TR U497 ( .A(n1344), .Y(n964) );
  CGENI_X1M_A9TR U498 ( .A(n1345), .B(n235), .CI(n820), .CON(n969) );
  INV_X0P7M_A9TR U499 ( .A(n1349), .Y(n1041) );
  CGENI_X1M_A9TR U500 ( .A(n1350), .B(n240), .CI(n762), .CON(n1046) );
  INV_X0P7M_A9TR U501 ( .A(n1354), .Y(n1034) );
  CGENI_X1M_A9TR U502 ( .A(n1355), .B(n245), .CI(n767), .CON(n1039) );
  INV_X0P7M_A9TR U503 ( .A(n1319), .Y(n1048) );
  CGENI_X1M_A9TR U504 ( .A(n1320), .B(n208), .CI(n840), .CON(n1053) );
  INV_X0P7M_A9TR U505 ( .A(n1324), .Y(n957) );
  CGENI_X1M_A9TR U506 ( .A(n1325), .B(n213), .CI(n825), .CON(n962) );
  INV_X0P7M_A9TR U507 ( .A(n1329), .Y(n950) );
  CGENI_X1M_A9TR U508 ( .A(n1330), .B(n218), .CI(n830), .CON(n955) );
  INV_X0P7M_A9TR U509 ( .A(n1334), .Y(n943) );
  CGENI_X1M_A9TR U510 ( .A(n1335), .B(n223), .CI(n835), .CON(n948) );
  AO21A1AI2_X0P7M_A9TR U511 ( .A0(n799), .A1(n798), .B0(n797), .C0(n796), .Y(
        \DUT_SM13_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U512 ( .A0(n804), .A1(n803), .B0(n802), .C0(n801), .Y(
        \DUT_SM14_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U513 ( .A0(n809), .A1(n808), .B0(n807), .C0(n806), .Y(
        \DUT_SM15_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U514 ( .A0(n814), .A1(n813), .B0(n812), .C0(n811), .Y(
        \DUT_SM16_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U515 ( .A0(n776), .A1(n775), .B0(n774), .C0(n773), .Y(
        \DUT_SM9_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U516 ( .A0(n782), .A1(n781), .B0(n780), .C0(n779), .Y(
        \DUT_SM10_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U517 ( .A0(n787), .A1(n786), .B0(n785), .C0(n784), .Y(
        \DUT_SM11_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U518 ( .A0(n793), .A1(n792), .B0(n791), .C0(n790), .Y(
        \DUT_SM12_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U519 ( .A0(n819), .A1(n818), .B0(n817), .C0(n816), .Y(
        \DUT_SM5_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U520 ( .A0(n824), .A1(n823), .B0(n822), .C0(n821), .Y(
        \DUT_SM6_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U521 ( .A0(n766), .A1(n765), .B0(n764), .C0(n763), .Y(
        \DUT_SM7_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U522 ( .A0(n771), .A1(n770), .B0(n769), .C0(n768), .Y(
        \DUT_SM8_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U523 ( .A0(n845), .A1(n844), .B0(n843), .C0(n842), .Y(
        \DUT_SM1_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U524 ( .A0(n829), .A1(n828), .B0(n827), .C0(n826), .Y(
        \DUT_SM2_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U525 ( .A0(n834), .A1(n833), .B0(n832), .C0(n831), .Y(
        \DUT_SM3_adjuster/N14 ) );
  AO21A1AI2_X0P7M_A9TR U526 ( .A0(n839), .A1(n838), .B0(n837), .C0(n836), .Y(
        \DUT_SM4_adjuster/N14 ) );
  AO21B_X0P7M_A9TR U527 ( .A0(n1169), .A1(SM13_issue_width_10_cycle[0]), .B0N(
        n739), .Y(\DUT_SM13_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U528 ( .A0(n1382), .A1(n738), .B0(n851), .C0(n1000), 
        .Y(n739) );
  AO21B_X0P7M_A9TR U529 ( .A0(n1174), .A1(SM14_issue_width_10_cycle[0]), .B0N(
        n737), .Y(\DUT_SM14_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U530 ( .A0(n1387), .A1(n736), .B0(n935), .C0(n993), .Y(
        n737) );
  AO21B_X0P7M_A9TR U531 ( .A0(n1179), .A1(SM15_issue_width_10_cycle[0]), .B0N(
        n735), .Y(\DUT_SM15_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U532 ( .A0(n1392), .A1(n734), .B0(n929), .C0(n986), .Y(
        n735) );
  AO21B_X0P7M_A9TR U533 ( .A0(n1183), .A1(SM16_issue_width_10_cycle[0]), .B0N(
        n761), .Y(\DUT_SM16_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U534 ( .A0(n1397), .A1(n760), .B0(n941), .C0(n979), .Y(
        n761) );
  AO21B_X0P7M_A9TR U535 ( .A0(n1149), .A1(SM9_issue_width_10_cycle[0]), .B0N(
        n747), .Y(\DUT_SM9_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U536 ( .A0(n1362), .A1(n746), .B0(n875), .C0(n1028), 
        .Y(n747) );
  AO21B_X0P7M_A9TR U537 ( .A0(n1154), .A1(SM10_issue_width_10_cycle[0]), .B0N(
        n745), .Y(\DUT_SM10_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U538 ( .A0(n1240), .A1(n744), .B0(n869), .C0(n1021), 
        .Y(n745) );
  AO21B_X0P7M_A9TR U539 ( .A0(n1159), .A1(SM11_issue_width_10_cycle[0]), .B0N(
        n743), .Y(\DUT_SM11_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U540 ( .A0(n1372), .A1(n742), .B0(n863), .C0(n1014), 
        .Y(n743) );
  AO21B_X0P7M_A9TR U541 ( .A0(n1164), .A1(SM12_issue_width_10_cycle[0]), .B0N(
        n741), .Y(\DUT_SM12_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U542 ( .A0(n1242), .A1(n740), .B0(n857), .C0(n1007), 
        .Y(n741) );
  AO21B_X0P7M_A9TR U543 ( .A0(n1129), .A1(SM5_issue_width_10_cycle[0]), .B0N(
        n755), .Y(\DUT_SM5_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U544 ( .A0(n1243), .A1(n754), .B0(n899), .C0(n972), .Y(
        n755) );
  AO21B_X0P7M_A9TR U545 ( .A0(n1134), .A1(SM6_issue_width_10_cycle[0]), .B0N(
        n753), .Y(\DUT_SM6_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U546 ( .A0(n1347), .A1(n752), .B0(n893), .C0(n965), .Y(
        n753) );
  AO21B_X0P7M_A9TR U547 ( .A0(n1139), .A1(SM7_issue_width_10_cycle[0]), .B0N(
        n751), .Y(\DUT_SM7_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U548 ( .A0(n1352), .A1(n750), .B0(n887), .C0(n1042), 
        .Y(n751) );
  AO21B_X0P7M_A9TR U549 ( .A0(n1144), .A1(SM8_issue_width_10_cycle[0]), .B0N(
        n749), .Y(\DUT_SM8_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U550 ( .A0(n1357), .A1(n748), .B0(n881), .C0(n1035), 
        .Y(n749) );
  AO21B_X0P7M_A9TR U551 ( .A0(n1109), .A1(SM1_issue_width_10_cycle[0]), .B0N(
        n733), .Y(\DUT_SM1_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U552 ( .A0(n1322), .A1(n732), .B0(n923), .C0(n1049), 
        .Y(n733) );
  AO21B_X0P7M_A9TR U553 ( .A0(n1114), .A1(SM2_issue_width_10_cycle[0]), .B0N(
        n731), .Y(\DUT_SM2_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U554 ( .A0(n1327), .A1(n730), .B0(n917), .C0(n958), .Y(
        n731) );
  AO21B_X0P7M_A9TR U555 ( .A0(n1119), .A1(SM3_issue_width_10_cycle[0]), .B0N(
        n759), .Y(\DUT_SM3_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U556 ( .A0(n1332), .A1(n758), .B0(n911), .C0(n951), .Y(
        n759) );
  AO21B_X0P7M_A9TR U557 ( .A0(n1124), .A1(SM4_issue_width_10_cycle[0]), .B0N(
        n757), .Y(\DUT_SM4_adjuster/N12 ) );
  AO21A1AI2_X0P7M_A9TR U558 ( .A0(n1337), .A1(n756), .B0(n905), .C0(n944), .Y(
        n757) );
  AO21A1AI2_X0P7M_A9TR U559 ( .A0(n851), .A1(n850), .B0(n849), .C0(n848), .Y(
        \DUT_SM13_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U560 ( .A0(n935), .A1(n934), .B0(n933), .C0(n932), .Y(
        \DUT_SM14_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U561 ( .A0(n929), .A1(n928), .B0(n927), .C0(n926), .Y(
        \DUT_SM15_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U562 ( .A0(n941), .A1(n940), .B0(n939), .C0(n938), .Y(
        \DUT_SM16_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U563 ( .A0(n875), .A1(n874), .B0(n873), .C0(n872), .Y(
        \DUT_SM9_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U564 ( .A0(n869), .A1(n868), .B0(n867), .C0(n866), .Y(
        \DUT_SM10_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U565 ( .A0(n863), .A1(n862), .B0(n861), .C0(n860), .Y(
        \DUT_SM11_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U566 ( .A0(n857), .A1(n856), .B0(n855), .C0(n854), .Y(
        \DUT_SM12_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U567 ( .A0(n899), .A1(n898), .B0(n897), .C0(n896), .Y(
        \DUT_SM5_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U568 ( .A0(n893), .A1(n892), .B0(n891), .C0(n890), .Y(
        \DUT_SM6_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U569 ( .A0(n887), .A1(n886), .B0(n885), .C0(n884), .Y(
        \DUT_SM7_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U570 ( .A0(n881), .A1(n880), .B0(n879), .C0(n878), .Y(
        \DUT_SM8_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U571 ( .A0(n923), .A1(n922), .B0(n921), .C0(n920), .Y(
        \DUT_SM1_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U572 ( .A0(n917), .A1(n916), .B0(n915), .C0(n914), .Y(
        \DUT_SM2_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U573 ( .A0(n911), .A1(n910), .B0(n909), .C0(n908), .Y(
        \DUT_SM3_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U574 ( .A0(n905), .A1(n904), .B0(n903), .C0(n902), .Y(
        \DUT_SM4_adjuster/N13 ) );
  AO21A1AI2_X0P7M_A9TR U575 ( .A0(n1004), .A1(n1003), .B0(n1002), .C0(n1001), 
        .Y(\DUT_SM13_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U576 ( .A0(n997), .A1(n996), .B0(n995), .C0(n994), .Y(
        \DUT_SM14_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U577 ( .A0(n990), .A1(n989), .B0(n988), .C0(n987), .Y(
        \DUT_SM15_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U578 ( .A0(n983), .A1(n982), .B0(n981), .C0(n980), .Y(
        \DUT_SM16_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U579 ( .A0(n1032), .A1(n1031), .B0(n1030), .C0(n1029), 
        .Y(\DUT_SM9_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U580 ( .A0(n1025), .A1(n1024), .B0(n1023), .C0(n1022), 
        .Y(\DUT_SM10_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U581 ( .A0(n1018), .A1(n1017), .B0(n1016), .C0(n1015), 
        .Y(\DUT_SM11_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U582 ( .A0(n1011), .A1(n1010), .B0(n1009), .C0(n1008), 
        .Y(\DUT_SM12_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U583 ( .A0(n976), .A1(n975), .B0(n974), .C0(n973), .Y(
        \DUT_SM5_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U584 ( .A0(n969), .A1(n968), .B0(n967), .C0(n966), .Y(
        \DUT_SM6_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U585 ( .A0(n1046), .A1(n1045), .B0(n1044), .C0(n1043), 
        .Y(\DUT_SM7_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U586 ( .A0(n1039), .A1(n1038), .B0(n1037), .C0(n1036), 
        .Y(\DUT_SM8_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U587 ( .A0(n1053), .A1(n1052), .B0(n1051), .C0(n1050), 
        .Y(\DUT_SM1_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U588 ( .A0(n962), .A1(n961), .B0(n960), .C0(n959), .Y(
        \DUT_SM2_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U589 ( .A0(n955), .A1(n954), .B0(n953), .C0(n952), .Y(
        \DUT_SM3_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U590 ( .A0(n948), .A1(n947), .B0(n946), .C0(n945), .Y(
        \DUT_SM4_adjuster/N15 ) );
  AO21A1AI2_X0P7M_A9TR U591 ( .A0(n277), .A1(SM13_issued_this_cycle[4]), .B0(
        n276), .C0(n275), .Y(\DUT_SM13_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U592 ( .A0(n282), .A1(SM14_issued_this_cycle[4]), .B0(
        n281), .C0(n280), .Y(\DUT_SM14_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U593 ( .A0(n287), .A1(SM15_issued_this_cycle[4]), .B0(
        n286), .C0(n285), .Y(\DUT_SM15_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U594 ( .A0(n293), .A1(SM16_issued_this_cycle[4]), .B0(
        n292), .C0(n291), .Y(\DUT_SM16_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U595 ( .A0(n255), .A1(SM9_issued_this_cycle[4]), .B0(
        n254), .C0(n253), .Y(\DUT_SM9_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U596 ( .A0(n261), .A1(SM10_issued_this_cycle[4]), .B0(
        n260), .C0(n259), .Y(\DUT_SM10_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U597 ( .A0(n266), .A1(SM11_issued_this_cycle[4]), .B0(
        n265), .C0(n264), .Y(\DUT_SM11_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U598 ( .A0(n272), .A1(SM12_issued_this_cycle[4]), .B0(
        n271), .C0(n270), .Y(\DUT_SM12_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U599 ( .A0(n234), .A1(SM5_issued_this_cycle[4]), .B0(
        n233), .C0(n232), .Y(\DUT_SM5_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U600 ( .A0(n239), .A1(SM6_issued_this_cycle[4]), .B0(
        n238), .C0(n237), .Y(\DUT_SM6_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U601 ( .A0(n244), .A1(SM7_issued_this_cycle[4]), .B0(
        n243), .C0(n242), .Y(\DUT_SM7_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U602 ( .A0(n249), .A1(SM8_issued_this_cycle[4]), .B0(
        n248), .C0(n247), .Y(\DUT_SM8_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U603 ( .A0(n212), .A1(SM1_issued_this_cycle[4]), .B0(
        n211), .C0(n210), .Y(\DUT_SM1_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U604 ( .A0(n217), .A1(SM2_issued_this_cycle[4]), .B0(
        n216), .C0(n215), .Y(\DUT_SM2_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U605 ( .A0(n222), .A1(SM3_issued_this_cycle[4]), .B0(
        n221), .C0(n220), .Y(\DUT_SM3_adjuster/N16 ) );
  AO21A1AI2_X0P7M_A9TR U606 ( .A0(n227), .A1(SM4_issued_this_cycle[4]), .B0(
        n226), .C0(n225), .Y(\DUT_SM4_adjuster/N16 ) );
  BUF_X5M_A9TR U607 ( .A(clk_controller), .Y(n1317) );
  BUFH_X11M_A9TR U608 ( .A(n1385), .Y(SM14_remaining[2]) );
  BUFH_X11M_A9TR U609 ( .A(n1390), .Y(SM15_remaining[2]) );
  BUFH_X11M_A9TR U610 ( .A(n1395), .Y(SM16_remaining[2]) );
  BUFH_X11M_A9TR U611 ( .A(n1360), .Y(SM9_remaining[2]) );
  BUFH_X11M_A9TR U612 ( .A(n1370), .Y(SM11_remaining[2]) );
  BUFH_X11M_A9TR U613 ( .A(n1340), .Y(SM5_remaining[2]) );
  BUFH_X11M_A9TR U614 ( .A(n1345), .Y(SM6_remaining[2]) );
  BUFH_X11M_A9TR U615 ( .A(n1350), .Y(SM7_remaining[2]) );
  BUFH_X11M_A9TR U616 ( .A(n1355), .Y(SM8_remaining[2]) );
  BUFH_X11M_A9TR U617 ( .A(n1325), .Y(SM2_remaining[2]) );
  BUFH_X11M_A9TR U618 ( .A(n1330), .Y(SM3_remaining[2]) );
  BUFH_X11M_A9TR U619 ( .A(n1335), .Y(SM4_remaining[2]) );
  BUFH_X11M_A9TR U620 ( .A(n1382), .Y(SM13_remaining[0]) );
  BUFH_X11M_A9TR U621 ( .A(n1387), .Y(SM14_remaining[0]) );
  BUFH_X11M_A9TR U622 ( .A(n1392), .Y(SM15_remaining[0]) );
  BUFH_X11M_A9TR U623 ( .A(n1397), .Y(SM16_remaining[0]) );
  BUFH_X11M_A9TR U624 ( .A(n1362), .Y(SM9_remaining[0]) );
  BUFH_X11M_A9TR U625 ( .A(n1372), .Y(SM11_remaining[0]) );
  BUFH_X11M_A9TR U626 ( .A(n1347), .Y(SM6_remaining[0]) );
  BUFH_X11M_A9TR U627 ( .A(n1352), .Y(SM7_remaining[0]) );
  BUFH_X11M_A9TR U628 ( .A(n1357), .Y(SM8_remaining[0]) );
  BUFH_X11M_A9TR U629 ( .A(n1322), .Y(SM1_remaining[0]) );
  BUFH_X11M_A9TR U630 ( .A(n1327), .Y(SM2_remaining[0]) );
  BUFH_X11M_A9TR U631 ( .A(n1332), .Y(SM3_remaining[0]) );
  BUFH_X11M_A9TR U632 ( .A(n1337), .Y(SM4_remaining[0]) );
  BUFH_X11M_A9TR U633 ( .A(n1318), .Y(SM1_remaining[4]) );
  INV_X0P7M_A9TR U634 ( .A(SM1_issued_this_cycle[2]), .Y(n208) );
  INV_X0P7M_A9TR U635 ( .A(SM1_issued_this_cycle[0]), .Y(n732) );
  CGENI_X1M_A9TR U636 ( .A(SM1_issued_this_cycle[1]), .B(n923), .CI(n919), 
        .CON(n840) );
  CGENI_X1M_A9TR U637 ( .A(n1053), .B(SM1_issued_this_cycle[3]), .CI(n1048), 
        .CON(n209) );
  XNOR2_X0P7M_A9TR U638 ( .A(n209), .B(n1318), .Y(n212) );
  BUFH_X1M_A9TR U639 ( .A(\DUT_SM16_adjuster/rst [0]), .Y(n1102) );
  INV_X0P7M_A9TR U640 ( .A(\DUT_SM1_adjuster/rst [2]), .Y(n1107) );
  NAND4BB_X0P5M_A9TR U641 ( .AN(\DUT_SM1_adjuster/rst [1]), .BN(
        \DUT_SM1_adjuster/rst [3]), .C(n1102), .D(n1107), .Y(n1049) );
  OAI21_X1M_A9TR U642 ( .A0(SM1_issued_this_cycle[4]), .A1(n212), .B0(n1049), 
        .Y(n211) );
  INV_X0P7M_A9TR U643 ( .A(n1049), .Y(n1109) );
  NAND2_X0P5A_A9TR U644 ( .A(n1109), .B(SM1_issue_width_10_cycle[4]), .Y(n210)
         );
  BUFH_X11M_A9TR U645 ( .A(n1323), .Y(SM2_remaining[4]) );
  INV_X0P7M_A9TR U646 ( .A(SM2_issued_this_cycle[2]), .Y(n213) );
  INV_X0P7M_A9TR U647 ( .A(SM2_issued_this_cycle[0]), .Y(n730) );
  CGENI_X1M_A9TR U648 ( .A(SM2_issued_this_cycle[1]), .B(n917), .CI(n913), 
        .CON(n825) );
  CGENI_X1M_A9TR U649 ( .A(n962), .B(SM2_issued_this_cycle[3]), .CI(n957), 
        .CON(n214) );
  XNOR2_X0P7M_A9TR U650 ( .A(n214), .B(n1323), .Y(n217) );
  INV_X0P7M_A9TR U651 ( .A(n1102), .Y(n1315) );
  INV_X0P7M_A9TR U652 ( .A(\DUT_SM2_adjuster/rst [2]), .Y(n1112) );
  NAND4BB_X0P5M_A9TR U653 ( .AN(\DUT_SM2_adjuster/rst [1]), .BN(
        \DUT_SM2_adjuster/rst [3]), .C(\DUT_SM16_adjuster/rst [0]), .D(n1112), 
        .Y(n958) );
  OAI21_X1M_A9TR U654 ( .A0(SM2_issued_this_cycle[4]), .A1(n217), .B0(n958), 
        .Y(n216) );
  INV_X0P7M_A9TR U655 ( .A(n958), .Y(n1114) );
  NAND2_X0P5A_A9TR U656 ( .A(n1114), .B(SM2_issue_width_10_cycle[4]), .Y(n215)
         );
  BUFH_X11M_A9TR U657 ( .A(n1328), .Y(SM3_remaining[4]) );
  INV_X0P7M_A9TR U658 ( .A(SM3_issued_this_cycle[2]), .Y(n218) );
  INV_X0P7M_A9TR U659 ( .A(SM3_issued_this_cycle[0]), .Y(n758) );
  CGENI_X1M_A9TR U660 ( .A(SM3_issued_this_cycle[1]), .B(n911), .CI(n907), 
        .CON(n830) );
  CGENI_X1M_A9TR U661 ( .A(n955), .B(SM3_issued_this_cycle[3]), .CI(n950), 
        .CON(n219) );
  XNOR2_X0P7M_A9TR U662 ( .A(n219), .B(n1328), .Y(n222) );
  INV_X0P7M_A9TR U663 ( .A(\DUT_SM3_adjuster/rst [2]), .Y(n1117) );
  NAND4BB_X0P5M_A9TR U664 ( .AN(\DUT_SM3_adjuster/rst [1]), .BN(
        \DUT_SM3_adjuster/rst [3]), .C(\DUT_SM16_adjuster/rst [0]), .D(n1117), 
        .Y(n951) );
  OAI21_X1M_A9TR U665 ( .A0(SM3_issued_this_cycle[4]), .A1(n222), .B0(n951), 
        .Y(n221) );
  INV_X0P7M_A9TR U666 ( .A(n951), .Y(n1119) );
  NAND2_X0P5A_A9TR U667 ( .A(n1119), .B(SM3_issue_width_10_cycle[4]), .Y(n220)
         );
  BUFH_X11M_A9TR U668 ( .A(n1333), .Y(SM4_remaining[4]) );
  INV_X0P7M_A9TR U669 ( .A(SM4_issued_this_cycle[2]), .Y(n223) );
  INV_X0P7M_A9TR U670 ( .A(SM4_issued_this_cycle[0]), .Y(n756) );
  CGENI_X1M_A9TR U671 ( .A(SM4_issued_this_cycle[1]), .B(n905), .CI(n901), 
        .CON(n835) );
  CGENI_X1M_A9TR U672 ( .A(n948), .B(SM4_issued_this_cycle[3]), .CI(n943), 
        .CON(n224) );
  XNOR2_X0P7M_A9TR U673 ( .A(n224), .B(n1333), .Y(n227) );
  INV_X0P7M_A9TR U674 ( .A(\DUT_SM4_adjuster/rst [2]), .Y(n1122) );
  NAND4BB_X0P5M_A9TR U675 ( .AN(\DUT_SM4_adjuster/rst [1]), .BN(
        \DUT_SM4_adjuster/rst [3]), .C(\DUT_SM16_adjuster/rst [0]), .D(n1122), 
        .Y(n944) );
  OAI21_X1M_A9TR U676 ( .A0(SM4_issued_this_cycle[4]), .A1(n227), .B0(n944), 
        .Y(n226) );
  INV_X0P7M_A9TR U677 ( .A(n944), .Y(n1124) );
  NAND2_X0P5A_A9TR U678 ( .A(n1124), .B(SM4_issue_width_10_cycle[4]), .Y(n225)
         );
  BUFH_X11M_A9TR U679 ( .A(n1338), .Y(SM5_remaining[4]) );
  BUFH_X1M_A9TR U680 ( .A(n1340), .Y(n230) );
  INV_X0P7M_A9TR U681 ( .A(SM5_issued_this_cycle[2]), .Y(n229) );
  INV_X0P7M_A9TR U682 ( .A(SM5_issued_this_cycle[0]), .Y(n754) );
  BUFH_X1M_A9TR U683 ( .A(n1342), .Y(n228) );
  CGENI_X1M_A9TR U684 ( .A(SM5_issued_this_cycle[1]), .B(n899), .CI(n895), 
        .CON(n815) );
  CGENI_X1M_A9TR U685 ( .A(n976), .B(SM5_issued_this_cycle[3]), .CI(n971), 
        .CON(n231) );
  XNOR2_X0P7M_A9TR U686 ( .A(n231), .B(n1338), .Y(n234) );
  INV_X0P7M_A9TR U687 ( .A(\DUT_SM5_adjuster/rst [2]), .Y(n1127) );
  NAND4BB_X0P5M_A9TR U688 ( .AN(\DUT_SM5_adjuster/rst [1]), .BN(
        \DUT_SM5_adjuster/rst [3]), .C(n1102), .D(n1127), .Y(n972) );
  OAI21_X1M_A9TR U689 ( .A0(SM5_issued_this_cycle[4]), .A1(n234), .B0(n972), 
        .Y(n233) );
  INV_X0P7M_A9TR U690 ( .A(n972), .Y(n1129) );
  NAND2_X0P5A_A9TR U691 ( .A(n1129), .B(SM5_issue_width_10_cycle[4]), .Y(n232)
         );
  BUFH_X11M_A9TR U692 ( .A(n1343), .Y(SM6_remaining[4]) );
  INV_X0P7M_A9TR U693 ( .A(SM6_issued_this_cycle[2]), .Y(n235) );
  INV_X0P7M_A9TR U694 ( .A(SM6_issued_this_cycle[0]), .Y(n752) );
  CGENI_X1M_A9TR U695 ( .A(SM6_issued_this_cycle[1]), .B(n893), .CI(n889), 
        .CON(n820) );
  CGENI_X1M_A9TR U696 ( .A(n969), .B(SM6_issued_this_cycle[3]), .CI(n964), 
        .CON(n236) );
  XNOR2_X0P7M_A9TR U697 ( .A(n236), .B(n1343), .Y(n239) );
  INV_X0P7M_A9TR U698 ( .A(\DUT_SM6_adjuster/rst [2]), .Y(n1132) );
  NAND4BB_X0P5M_A9TR U699 ( .AN(\DUT_SM6_adjuster/rst [1]), .BN(
        \DUT_SM6_adjuster/rst [3]), .C(\DUT_SM16_adjuster/rst [0]), .D(n1132), 
        .Y(n965) );
  OAI21_X1M_A9TR U700 ( .A0(SM6_issued_this_cycle[4]), .A1(n239), .B0(n965), 
        .Y(n238) );
  INV_X0P7M_A9TR U701 ( .A(n965), .Y(n1134) );
  NAND2_X0P5A_A9TR U702 ( .A(n1134), .B(SM6_issue_width_10_cycle[4]), .Y(n237)
         );
  BUFH_X11M_A9TR U703 ( .A(n1348), .Y(SM7_remaining[4]) );
  INV_X0P7M_A9TR U704 ( .A(SM7_issued_this_cycle[2]), .Y(n240) );
  INV_X0P7M_A9TR U705 ( .A(SM7_issued_this_cycle[0]), .Y(n750) );
  CGENI_X1M_A9TR U706 ( .A(SM7_issued_this_cycle[1]), .B(n887), .CI(n883), 
        .CON(n762) );
  CGENI_X1M_A9TR U707 ( .A(n1046), .B(SM7_issued_this_cycle[3]), .CI(n1041), 
        .CON(n241) );
  XNOR2_X0P7M_A9TR U708 ( .A(n241), .B(n1348), .Y(n244) );
  INV_X0P7M_A9TR U709 ( .A(\DUT_SM7_adjuster/rst [2]), .Y(n1137) );
  NAND4BB_X0P5M_A9TR U710 ( .AN(\DUT_SM7_adjuster/rst [1]), .BN(
        \DUT_SM7_adjuster/rst [3]), .C(n1102), .D(n1137), .Y(n1042) );
  OAI21_X1M_A9TR U711 ( .A0(SM7_issued_this_cycle[4]), .A1(n244), .B0(n1042), 
        .Y(n243) );
  INV_X0P7M_A9TR U712 ( .A(n1042), .Y(n1139) );
  NAND2_X0P5A_A9TR U713 ( .A(n1139), .B(SM7_issue_width_10_cycle[4]), .Y(n242)
         );
  BUFH_X11M_A9TR U714 ( .A(n1353), .Y(SM8_remaining[4]) );
  INV_X0P7M_A9TR U715 ( .A(SM8_issued_this_cycle[2]), .Y(n245) );
  INV_X0P7M_A9TR U716 ( .A(SM8_issued_this_cycle[0]), .Y(n748) );
  CGENI_X1M_A9TR U717 ( .A(SM8_issued_this_cycle[1]), .B(n881), .CI(n877), 
        .CON(n767) );
  CGENI_X1M_A9TR U718 ( .A(n1039), .B(SM8_issued_this_cycle[3]), .CI(n1034), 
        .CON(n246) );
  XNOR2_X0P7M_A9TR U719 ( .A(n246), .B(n1353), .Y(n249) );
  INV_X0P7M_A9TR U720 ( .A(\DUT_SM8_adjuster/rst [2]), .Y(n1142) );
  NAND4BB_X0P5M_A9TR U721 ( .AN(\DUT_SM8_adjuster/rst [1]), .BN(
        \DUT_SM8_adjuster/rst [3]), .C(n1102), .D(n1142), .Y(n1035) );
  OAI21_X1M_A9TR U722 ( .A0(SM8_issued_this_cycle[4]), .A1(n249), .B0(n1035), 
        .Y(n248) );
  INV_X0P7M_A9TR U723 ( .A(n1035), .Y(n1144) );
  NAND2_X0P5A_A9TR U724 ( .A(n1144), .B(SM8_issue_width_10_cycle[4]), .Y(n247)
         );
  BUFH_X11M_A9TR U725 ( .A(n1358), .Y(SM9_remaining[4]) );
  BUFH_X1M_A9TR U726 ( .A(n1360), .Y(n251) );
  INV_X0P7M_A9TR U727 ( .A(SM9_issued_this_cycle[2]), .Y(n250) );
  INV_X0P7M_A9TR U728 ( .A(SM9_issued_this_cycle[0]), .Y(n746) );
  CGENI_X1M_A9TR U729 ( .A(SM9_issued_this_cycle[1]), .B(n875), .CI(n871), 
        .CON(n772) );
  CGENI_X1M_A9TR U730 ( .A(n1032), .B(SM9_issued_this_cycle[3]), .CI(n1027), 
        .CON(n252) );
  XNOR2_X0P7M_A9TR U731 ( .A(n252), .B(n1358), .Y(n255) );
  INV_X0P7M_A9TR U732 ( .A(\DUT_SM9_adjuster/rst [2]), .Y(n1147) );
  NAND4BB_X0P5M_A9TR U733 ( .AN(\DUT_SM9_adjuster/rst [1]), .BN(
        \DUT_SM9_adjuster/rst [3]), .C(n1102), .D(n1147), .Y(n1028) );
  OAI21_X1M_A9TR U734 ( .A0(SM9_issued_this_cycle[4]), .A1(n255), .B0(n1028), 
        .Y(n254) );
  INV_X0P7M_A9TR U735 ( .A(n1028), .Y(n1149) );
  NAND2_X0P5A_A9TR U736 ( .A(n1149), .B(SM9_issue_width_10_cycle[4]), .Y(n253)
         );
  BUFH_X11M_A9TR U737 ( .A(n1363), .Y(SM10_remaining[4]) );
  INV_X0P7M_A9TR U738 ( .A(SM10_issued_this_cycle[2]), .Y(n257) );
  INV_X0P7M_A9TR U739 ( .A(SM10_issued_this_cycle[0]), .Y(n744) );
  BUFH_X1M_A9TR U740 ( .A(n1367), .Y(n256) );
  CGENI_X1M_A9TR U741 ( .A(SM10_issued_this_cycle[1]), .B(n869), .CI(n865), 
        .CON(n777) );
  CGENI_X1M_A9TR U742 ( .A(n1025), .B(SM10_issued_this_cycle[3]), .CI(n1020), 
        .CON(n258) );
  XNOR2_X0P7M_A9TR U743 ( .A(n258), .B(n1363), .Y(n261) );
  INV_X0P7M_A9TR U744 ( .A(\DUT_SM10_adjuster/rst [2]), .Y(n1152) );
  NAND4BB_X0P5M_A9TR U745 ( .AN(\DUT_SM10_adjuster/rst [1]), .BN(
        \DUT_SM10_adjuster/rst [3]), .C(n1102), .D(n1152), .Y(n1021) );
  OAI21_X1M_A9TR U746 ( .A0(SM10_issued_this_cycle[4]), .A1(n261), .B0(n1021), 
        .Y(n260) );
  INV_X0P7M_A9TR U747 ( .A(n1021), .Y(n1154) );
  NAND2_X0P5A_A9TR U748 ( .A(n1154), .B(SM10_issue_width_10_cycle[4]), .Y(n259) );
  BUFH_X11M_A9TR U749 ( .A(n1368), .Y(SM11_remaining[4]) );
  INV_X0P7M_A9TR U750 ( .A(SM11_issued_this_cycle[2]), .Y(n262) );
  INV_X0P7M_A9TR U751 ( .A(SM11_issued_this_cycle[0]), .Y(n742) );
  CGENI_X1M_A9TR U752 ( .A(SM11_issued_this_cycle[1]), .B(n863), .CI(n859), 
        .CON(n783) );
  CGENI_X1M_A9TR U753 ( .A(n1018), .B(SM11_issued_this_cycle[3]), .CI(n1013), 
        .CON(n263) );
  XNOR2_X0P7M_A9TR U754 ( .A(n263), .B(n1368), .Y(n266) );
  INV_X0P7M_A9TR U755 ( .A(\DUT_SM11_adjuster/rst [2]), .Y(n1157) );
  NAND4BB_X0P5M_A9TR U756 ( .AN(\DUT_SM11_adjuster/rst [1]), .BN(
        \DUT_SM11_adjuster/rst [3]), .C(n1102), .D(n1157), .Y(n1014) );
  OAI21_X1M_A9TR U757 ( .A0(SM11_issued_this_cycle[4]), .A1(n266), .B0(n1014), 
        .Y(n265) );
  INV_X0P7M_A9TR U758 ( .A(n1014), .Y(n1159) );
  NAND2_X0P5A_A9TR U759 ( .A(n1159), .B(SM11_issue_width_10_cycle[4]), .Y(n264) );
  BUFH_X11M_A9TR U760 ( .A(n1373), .Y(SM12_remaining[4]) );
  INV_X0P7M_A9TR U761 ( .A(SM12_issued_this_cycle[2]), .Y(n268) );
  INV_X0P7M_A9TR U762 ( .A(SM12_issued_this_cycle[0]), .Y(n740) );
  BUFH_X1M_A9TR U763 ( .A(n1377), .Y(n267) );
  CGENI_X1M_A9TR U764 ( .A(SM12_issued_this_cycle[1]), .B(n857), .CI(n853), 
        .CON(n788) );
  CGENI_X1M_A9TR U765 ( .A(n1011), .B(SM12_issued_this_cycle[3]), .CI(n1006), 
        .CON(n269) );
  XNOR2_X0P7M_A9TR U766 ( .A(n269), .B(n1373), .Y(n272) );
  INV_X0P7M_A9TR U767 ( .A(\DUT_SM12_adjuster/rst [2]), .Y(n1162) );
  NAND4BB_X0P5M_A9TR U768 ( .AN(\DUT_SM12_adjuster/rst [1]), .BN(
        \DUT_SM12_adjuster/rst [3]), .C(n1102), .D(n1162), .Y(n1007) );
  OAI21_X1M_A9TR U769 ( .A0(SM12_issued_this_cycle[4]), .A1(n272), .B0(n1007), 
        .Y(n271) );
  INV_X0P7M_A9TR U770 ( .A(n1007), .Y(n1164) );
  NAND2_X0P5A_A9TR U771 ( .A(n1164), .B(SM12_issue_width_10_cycle[4]), .Y(n270) );
  BUFH_X11M_A9TR U772 ( .A(n1378), .Y(SM13_remaining[4]) );
  INV_X0P7M_A9TR U773 ( .A(SM13_issued_this_cycle[2]), .Y(n273) );
  INV_X0P7M_A9TR U774 ( .A(SM13_issued_this_cycle[0]), .Y(n738) );
  CGENI_X1M_A9TR U775 ( .A(SM13_issued_this_cycle[1]), .B(n851), .CI(n847), 
        .CON(n794) );
  CGENI_X1M_A9TR U776 ( .A(n1004), .B(SM13_issued_this_cycle[3]), .CI(n999), 
        .CON(n274) );
  XNOR2_X0P7M_A9TR U777 ( .A(n274), .B(n1378), .Y(n277) );
  INV_X0P7M_A9TR U778 ( .A(\DUT_SM13_adjuster/rst [2]), .Y(n1167) );
  NAND4BB_X0P5M_A9TR U779 ( .AN(\DUT_SM13_adjuster/rst [1]), .BN(
        \DUT_SM13_adjuster/rst [3]), .C(n1102), .D(n1167), .Y(n1000) );
  OAI21_X1M_A9TR U780 ( .A0(SM13_issued_this_cycle[4]), .A1(n277), .B0(n1000), 
        .Y(n276) );
  INV_X0P7M_A9TR U781 ( .A(n1000), .Y(n1169) );
  NAND2_X0P5A_A9TR U782 ( .A(n1169), .B(SM13_issue_width_10_cycle[4]), .Y(n275) );
  BUFH_X11M_A9TR U783 ( .A(n1383), .Y(SM14_remaining[4]) );
  INV_X0P7M_A9TR U784 ( .A(SM14_issued_this_cycle[2]), .Y(n278) );
  INV_X0P7M_A9TR U785 ( .A(SM14_issued_this_cycle[0]), .Y(n736) );
  CGENI_X1M_A9TR U786 ( .A(SM14_issued_this_cycle[1]), .B(n935), .CI(n931), 
        .CON(n800) );
  CGENI_X1M_A9TR U787 ( .A(n997), .B(SM14_issued_this_cycle[3]), .CI(n992), 
        .CON(n279) );
  XNOR2_X0P7M_A9TR U788 ( .A(n279), .B(n1383), .Y(n282) );
  INV_X0P7M_A9TR U789 ( .A(\DUT_SM14_adjuster/rst [2]), .Y(n1172) );
  NAND4BB_X0P5M_A9TR U790 ( .AN(\DUT_SM14_adjuster/rst [1]), .BN(
        \DUT_SM14_adjuster/rst [3]), .C(n1102), .D(n1172), .Y(n993) );
  OAI21_X1M_A9TR U791 ( .A0(SM14_issued_this_cycle[4]), .A1(n282), .B0(n993), 
        .Y(n281) );
  INV_X0P7M_A9TR U792 ( .A(n993), .Y(n1174) );
  NAND2_X0P5A_A9TR U793 ( .A(n1174), .B(SM14_issue_width_10_cycle[4]), .Y(n280) );
  BUFH_X11M_A9TR U794 ( .A(n1388), .Y(SM15_remaining[4]) );
  INV_X0P7M_A9TR U795 ( .A(SM15_issued_this_cycle[2]), .Y(n283) );
  INV_X0P7M_A9TR U796 ( .A(SM15_issued_this_cycle[0]), .Y(n734) );
  CGENI_X1M_A9TR U797 ( .A(SM15_issued_this_cycle[1]), .B(n929), .CI(n925), 
        .CON(n805) );
  CGENI_X1M_A9TR U798 ( .A(n990), .B(SM15_issued_this_cycle[3]), .CI(n985), 
        .CON(n284) );
  XNOR2_X0P7M_A9TR U799 ( .A(n284), .B(n1388), .Y(n287) );
  INV_X0P7M_A9TR U800 ( .A(\DUT_SM15_adjuster/rst [2]), .Y(n1177) );
  NAND4BB_X0P5M_A9TR U801 ( .AN(\DUT_SM15_adjuster/rst [1]), .BN(
        \DUT_SM15_adjuster/rst [3]), .C(\DUT_SM16_adjuster/rst [0]), .D(n1177), 
        .Y(n986) );
  OAI21_X1M_A9TR U802 ( .A0(SM15_issued_this_cycle[4]), .A1(n287), .B0(n986), 
        .Y(n286) );
  INV_X0P7M_A9TR U803 ( .A(n986), .Y(n1179) );
  NAND2_X0P5A_A9TR U804 ( .A(n1179), .B(SM15_issue_width_10_cycle[4]), .Y(n285) );
  BUFH_X11M_A9TR U805 ( .A(n1393), .Y(SM16_remaining[4]) );
  BUFH_X1M_A9TR U806 ( .A(n1395), .Y(n289) );
  INV_X0P7M_A9TR U807 ( .A(SM16_issued_this_cycle[2]), .Y(n288) );
  INV_X0P7M_A9TR U808 ( .A(SM16_issued_this_cycle[0]), .Y(n760) );
  CGENI_X1M_A9TR U809 ( .A(SM16_issued_this_cycle[1]), .B(n941), .CI(n937), 
        .CON(n810) );
  CGENI_X1M_A9TR U810 ( .A(n983), .B(SM16_issued_this_cycle[3]), .CI(n978), 
        .CON(n290) );
  XNOR2_X0P7M_A9TR U811 ( .A(n290), .B(n1393), .Y(n293) );
  NAND4BB_X0P5M_A9TR U812 ( .AN(\DUT_SM16_adjuster/rst [1]), .BN(
        \DUT_SM16_adjuster/rst [3]), .C(n1102), .D(n1316), .Y(n979) );
  OAI21_X1M_A9TR U813 ( .A0(SM16_issued_this_cycle[4]), .A1(n293), .B0(n979), 
        .Y(n292) );
  INV_X0P7M_A9TR U814 ( .A(n979), .Y(n1183) );
  NAND2_X0P5A_A9TR U815 ( .A(n1183), .B(SM16_issue_width_10_cycle[4]), .Y(n291) );
  BUFH_X11M_A9TR U816 ( .A(n1319), .Y(SM1_remaining[3]) );
  BUFH_X11M_A9TR U817 ( .A(n1324), .Y(SM2_remaining[3]) );
  BUFH_X11M_A9TR U818 ( .A(n1329), .Y(SM3_remaining[3]) );
  BUFH_X11M_A9TR U819 ( .A(n1334), .Y(SM4_remaining[3]) );
  BUFH_X11M_A9TR U820 ( .A(n1339), .Y(SM5_remaining[3]) );
  BUFH_X11M_A9TR U821 ( .A(n1344), .Y(SM6_remaining[3]) );
  BUFH_X11M_A9TR U822 ( .A(n1349), .Y(SM7_remaining[3]) );
  BUFH_X11M_A9TR U823 ( .A(n1354), .Y(SM8_remaining[3]) );
  BUFH_X11M_A9TR U824 ( .A(n1359), .Y(SM9_remaining[3]) );
  BUFH_X11M_A9TR U825 ( .A(n1364), .Y(SM10_remaining[3]) );
  BUFH_X11M_A9TR U826 ( .A(n1369), .Y(SM11_remaining[3]) );
  BUFH_X11M_A9TR U827 ( .A(n1374), .Y(SM12_remaining[3]) );
  BUFH_X11M_A9TR U828 ( .A(n1379), .Y(SM13_remaining[3]) );
  BUFH_X11M_A9TR U829 ( .A(n1384), .Y(SM14_remaining[3]) );
  BUFH_X11M_A9TR U830 ( .A(n1389), .Y(SM15_remaining[3]) );
  BUFH_X11M_A9TR U831 ( .A(n1394), .Y(SM16_remaining[3]) );
  BUFH_X11M_A9TR U832 ( .A(n1321), .Y(SM1_remaining[1]) );
  BUFH_X11M_A9TR U833 ( .A(n1326), .Y(SM2_remaining[1]) );
  BUFH_X11M_A9TR U834 ( .A(n1331), .Y(SM3_remaining[1]) );
  BUFH_X11M_A9TR U835 ( .A(n1336), .Y(SM4_remaining[1]) );
  BUFH_X11M_A9TR U836 ( .A(n1341), .Y(SM5_remaining[1]) );
  BUFH_X11M_A9TR U837 ( .A(n1346), .Y(SM6_remaining[1]) );
  BUFH_X11M_A9TR U838 ( .A(n1351), .Y(SM7_remaining[1]) );
  BUFH_X11M_A9TR U839 ( .A(n1356), .Y(SM8_remaining[1]) );
  BUFH_X11M_A9TR U840 ( .A(n1361), .Y(SM9_remaining[1]) );
  BUFH_X11M_A9TR U841 ( .A(n1366), .Y(SM10_remaining[1]) );
  BUFH_X11M_A9TR U842 ( .A(n1371), .Y(SM11_remaining[1]) );
  BUFH_X11M_A9TR U843 ( .A(n1376), .Y(SM12_remaining[1]) );
  BUFH_X11M_A9TR U844 ( .A(n1381), .Y(SM13_remaining[1]) );
  BUFH_X11M_A9TR U845 ( .A(n1386), .Y(SM14_remaining[1]) );
  BUFH_X11M_A9TR U846 ( .A(n1391), .Y(SM15_remaining[1]) );
  BUFH_X11M_A9TR U847 ( .A(n1396), .Y(SM16_remaining[1]) );
  INV_X0P7M_A9TR U848 ( .A(SM8_voltage[7]), .Y(n295) );
  OAI21_X1M_A9TR U849 ( .A0(n295), .A1(SM8_voltage[5]), .B0(SM8_voltage[6]), 
        .Y(n297) );
  INV_X0P7M_A9TR U850 ( .A(n297), .Y(n303) );
  NOR3_X0P7A_A9TR U851 ( .A(SM8_voltage[5]), .B(SM8_voltage[6]), .C(n295), .Y(
        n296) );
  NOR2_X0P7A_A9TR U852 ( .A(n303), .B(n296), .Y(n302) );
  INV_X0P7M_A9TR U853 ( .A(SM8_voltage[4]), .Y(n298) );
  OAI21_X1M_A9TR U854 ( .A0(SM8_voltage[5]), .A1(SM8_voltage[6]), .B0(
        SM8_voltage[7]), .Y(n319) );
  NOR2_X0P7A_A9TR U855 ( .A(SM8_voltage[5]), .B(n319), .Y(n294) );
  AOI21_X0P7M_A9TR U856 ( .A0(SM8_voltage[5]), .A1(n295), .B0(n294), .Y(n301)
         );
  INV_X0P7M_A9TR U857 ( .A(n296), .Y(n299) );
  AO21A1AI2_X0P7M_A9TR U858 ( .A0(n298), .A1(n301), .B0(n297), .C0(n299), .Y(
        n1056) );
  NOR2B_X1M_A9TR U859 ( .AN(n1056), .B(SM8_voltage[4]), .Y(n300) );
  AOI21_X0P7M_A9TR U860 ( .A0(n302), .A1(SM8_voltage[4]), .B0(n300), .Y(n306)
         );
  NAND2B_X0P5M_A9TR U861 ( .AN(SM8_voltage[3]), .B(n306), .Y(n304) );
  OAI22_X0P5M_A9TR U862 ( .A0(n301), .A1(n300), .B0(SM8_voltage[4]), .B1(n299), 
        .Y(n310) );
  AOI21_X0P7M_A9TR U863 ( .A0(n303), .A1(n1056), .B0(n302), .Y(n308) );
  AOI21_X0P7M_A9TR U864 ( .A0(n304), .A1(n310), .B0(n308), .Y(n1212) );
  XNOR2_X0P7M_A9TR U865 ( .A(SM8_voltage[3]), .B(n1212), .Y(n313) );
  NOR2_X0P7A_A9TR U866 ( .A(SM8_voltage[3]), .B(n1212), .Y(n307) );
  NAND2_X0P5A_A9TR U867 ( .A(n306), .B(n308), .Y(n305) );
  OAI22_X0P5M_A9TR U868 ( .A0(n307), .A1(n306), .B0(n305), .B1(SM8_voltage[3]), 
        .Y(n317) );
  INV_X0P7M_A9TR U869 ( .A(n310), .Y(n309) );
  AOI22_X0P7M_A9TR U870 ( .A0(n310), .A1(n1212), .B0(n309), .B1(n308), .Y(n318) );
  INV_X0P7M_A9TR U871 ( .A(n318), .Y(n311) );
  OA21A1OI2_X0P5M_A9TR U872 ( .A0(SM8_voltage[2]), .A1(n313), .B0(n317), .C0(
        n311), .Y(n315) );
  INV_X0P7M_A9TR U873 ( .A(n315), .Y(n1054) );
  CGENI_X1M_A9TR U874 ( .A(n315), .B(SM8_voltage[1]), .CI(SM8_voltage[2]), 
        .CON(n312) );
  NOR2B_X1M_A9TR U875 ( .AN(n313), .B(n312), .Y(n314) );
  AOI21_X0P7M_A9TR U876 ( .A0(n315), .A1(n317), .B0(n314), .Y(n316) );
  OAI21_X1M_A9TR U877 ( .A0(n318), .A1(n317), .B0(n316), .Y(
        \DUT_controller/N75 ) );
  NOR2_X0P7A_A9TR U878 ( .A(n1054), .B(\DUT_controller/N75 ), .Y(n1213) );
  NOR2_X0P7A_A9TR U879 ( .A(n1212), .B(n1213), .Y(n1211) );
  NOR2_X0P7A_A9TR U880 ( .A(n1211), .B(n1056), .Y(n1055) );
  XNOR2_X0P7M_A9TR U881 ( .A(n1055), .B(n319), .Y(\DUT_controller/N79 ) );
  INV_X0P7M_A9TR U882 ( .A(SM16_voltage[7]), .Y(n321) );
  OAI21_X1M_A9TR U883 ( .A0(n321), .A1(SM16_voltage[5]), .B0(SM16_voltage[6]), 
        .Y(n323) );
  INV_X0P7M_A9TR U884 ( .A(n323), .Y(n329) );
  NOR3_X0P7A_A9TR U885 ( .A(SM16_voltage[5]), .B(SM16_voltage[6]), .C(n321), 
        .Y(n322) );
  NOR2_X0P7A_A9TR U886 ( .A(n329), .B(n322), .Y(n328) );
  INV_X0P7M_A9TR U887 ( .A(SM16_voltage[4]), .Y(n324) );
  OAI21_X1M_A9TR U888 ( .A0(SM16_voltage[5]), .A1(SM16_voltage[6]), .B0(
        SM16_voltage[7]), .Y(n345) );
  NOR2_X0P7A_A9TR U889 ( .A(SM16_voltage[5]), .B(n345), .Y(n320) );
  AOI21_X0P7M_A9TR U890 ( .A0(SM16_voltage[5]), .A1(n321), .B0(n320), .Y(n327)
         );
  INV_X0P7M_A9TR U891 ( .A(n322), .Y(n325) );
  AO21A1AI2_X0P7M_A9TR U892 ( .A0(n324), .A1(n327), .B0(n323), .C0(n325), .Y(
        n1062) );
  NOR2B_X1M_A9TR U893 ( .AN(n1062), .B(SM16_voltage[4]), .Y(n326) );
  AOI21_X0P7M_A9TR U894 ( .A0(n328), .A1(SM16_voltage[4]), .B0(n326), .Y(n332)
         );
  NAND2B_X0P5M_A9TR U895 ( .AN(SM16_voltage[3]), .B(n332), .Y(n330) );
  OAI22_X0P5M_A9TR U896 ( .A0(n327), .A1(n326), .B0(SM16_voltage[4]), .B1(n325), .Y(n336) );
  AOI21_X0P7M_A9TR U897 ( .A0(n329), .A1(n1062), .B0(n328), .Y(n334) );
  AOI21_X0P7M_A9TR U898 ( .A0(n330), .A1(n336), .B0(n334), .Y(n1188) );
  XNOR2_X0P7M_A9TR U899 ( .A(SM16_voltage[3]), .B(n1188), .Y(n339) );
  NOR2_X0P7A_A9TR U900 ( .A(SM16_voltage[3]), .B(n1188), .Y(n333) );
  NAND2_X0P5A_A9TR U901 ( .A(n332), .B(n334), .Y(n331) );
  OAI22_X0P5M_A9TR U902 ( .A0(n333), .A1(n332), .B0(n331), .B1(SM16_voltage[3]), .Y(n343) );
  INV_X0P7M_A9TR U903 ( .A(n336), .Y(n335) );
  AOI22_X0P7M_A9TR U904 ( .A0(n336), .A1(n1188), .B0(n335), .B1(n334), .Y(n344) );
  INV_X0P7M_A9TR U905 ( .A(n344), .Y(n337) );
  OA21A1OI2_X0P5M_A9TR U906 ( .A0(SM16_voltage[2]), .A1(n339), .B0(n343), .C0(
        n337), .Y(n341) );
  INV_X0P7M_A9TR U907 ( .A(n341), .Y(n1060) );
  CGENI_X1M_A9TR U908 ( .A(n341), .B(SM16_voltage[1]), .CI(SM16_voltage[2]), 
        .CON(n338) );
  NOR2B_X1M_A9TR U909 ( .AN(n339), .B(n338), .Y(n340) );
  AOI21_X0P7M_A9TR U910 ( .A0(n341), .A1(n343), .B0(n340), .Y(n342) );
  OAI21_X1M_A9TR U911 ( .A0(n344), .A1(n343), .B0(n342), .Y(
        \DUT_controller/N155 ) );
  NOR2_X0P7A_A9TR U912 ( .A(n1060), .B(\DUT_controller/N155 ), .Y(n1189) );
  NOR2_X0P7A_A9TR U913 ( .A(n1188), .B(n1189), .Y(n1187) );
  NOR2_X0P7A_A9TR U914 ( .A(n1187), .B(n1062), .Y(n1061) );
  XNOR2_X0P7M_A9TR U915 ( .A(n1061), .B(n345), .Y(\DUT_controller/N159 ) );
  INV_X0P7M_A9TR U916 ( .A(SM15_voltage[7]), .Y(n347) );
  OAI21_X1M_A9TR U917 ( .A0(n347), .A1(SM15_voltage[5]), .B0(SM15_voltage[6]), 
        .Y(n349) );
  INV_X0P7M_A9TR U918 ( .A(n349), .Y(n355) );
  NOR3_X0P7A_A9TR U919 ( .A(SM15_voltage[5]), .B(SM15_voltage[6]), .C(n347), 
        .Y(n348) );
  NOR2_X0P7A_A9TR U920 ( .A(n355), .B(n348), .Y(n354) );
  INV_X0P7M_A9TR U921 ( .A(SM15_voltage[4]), .Y(n350) );
  OAI21_X1M_A9TR U922 ( .A0(SM15_voltage[5]), .A1(SM15_voltage[6]), .B0(
        SM15_voltage[7]), .Y(n371) );
  NOR2_X0P7A_A9TR U923 ( .A(SM15_voltage[5]), .B(n371), .Y(n346) );
  AOI21_X0P7M_A9TR U924 ( .A0(SM15_voltage[5]), .A1(n347), .B0(n346), .Y(n353)
         );
  INV_X0P7M_A9TR U925 ( .A(n348), .Y(n351) );
  AO21A1AI2_X0P7M_A9TR U926 ( .A0(n350), .A1(n353), .B0(n349), .C0(n351), .Y(
        n1065) );
  NOR2B_X1M_A9TR U927 ( .AN(n1065), .B(SM15_voltage[4]), .Y(n352) );
  AOI21_X0P7M_A9TR U928 ( .A0(n354), .A1(SM15_voltage[4]), .B0(n352), .Y(n358)
         );
  NAND2B_X0P5M_A9TR U929 ( .AN(SM15_voltage[3]), .B(n358), .Y(n356) );
  OAI22_X0P5M_A9TR U930 ( .A0(n353), .A1(n352), .B0(SM15_voltage[4]), .B1(n351), .Y(n362) );
  AOI21_X0P7M_A9TR U931 ( .A0(n355), .A1(n1065), .B0(n354), .Y(n360) );
  AOI21_X0P7M_A9TR U932 ( .A0(n356), .A1(n362), .B0(n360), .Y(n1191) );
  XNOR2_X0P7M_A9TR U933 ( .A(SM15_voltage[3]), .B(n1191), .Y(n365) );
  NOR2_X0P7A_A9TR U934 ( .A(SM15_voltage[3]), .B(n1191), .Y(n359) );
  NAND2_X0P5A_A9TR U935 ( .A(n358), .B(n360), .Y(n357) );
  OAI22_X0P5M_A9TR U936 ( .A0(n359), .A1(n358), .B0(n357), .B1(SM15_voltage[3]), .Y(n369) );
  INV_X0P7M_A9TR U937 ( .A(n362), .Y(n361) );
  AOI22_X0P7M_A9TR U938 ( .A0(n362), .A1(n1191), .B0(n361), .B1(n360), .Y(n370) );
  INV_X0P7M_A9TR U939 ( .A(n370), .Y(n363) );
  OA21A1OI2_X0P5M_A9TR U940 ( .A0(SM15_voltage[2]), .A1(n365), .B0(n369), .C0(
        n363), .Y(n367) );
  INV_X0P7M_A9TR U941 ( .A(n367), .Y(n1063) );
  CGENI_X1M_A9TR U942 ( .A(n367), .B(SM15_voltage[1]), .CI(SM15_voltage[2]), 
        .CON(n364) );
  NOR2B_X1M_A9TR U943 ( .AN(n365), .B(n364), .Y(n366) );
  AOI21_X0P7M_A9TR U944 ( .A0(n367), .A1(n369), .B0(n366), .Y(n368) );
  OAI21_X1M_A9TR U945 ( .A0(n370), .A1(n369), .B0(n368), .Y(
        \DUT_controller/N145 ) );
  NOR2_X0P7A_A9TR U946 ( .A(n1063), .B(\DUT_controller/N145 ), .Y(n1192) );
  NOR2_X0P7A_A9TR U947 ( .A(n1191), .B(n1192), .Y(n1190) );
  NOR2_X0P7A_A9TR U948 ( .A(n1190), .B(n1065), .Y(n1064) );
  XNOR2_X0P7M_A9TR U949 ( .A(n1064), .B(n371), .Y(\DUT_controller/N149 ) );
  INV_X0P7M_A9TR U950 ( .A(SM14_voltage[7]), .Y(n373) );
  OAI21_X1M_A9TR U951 ( .A0(n373), .A1(SM14_voltage[5]), .B0(SM14_voltage[6]), 
        .Y(n375) );
  INV_X0P7M_A9TR U952 ( .A(n375), .Y(n381) );
  NOR3_X0P7A_A9TR U953 ( .A(SM14_voltage[5]), .B(SM14_voltage[6]), .C(n373), 
        .Y(n374) );
  NOR2_X0P7A_A9TR U954 ( .A(n381), .B(n374), .Y(n380) );
  INV_X0P7M_A9TR U955 ( .A(SM14_voltage[4]), .Y(n376) );
  OAI21_X1M_A9TR U956 ( .A0(SM14_voltage[5]), .A1(SM14_voltage[6]), .B0(
        SM14_voltage[7]), .Y(n397) );
  NOR2_X0P7A_A9TR U957 ( .A(SM14_voltage[5]), .B(n397), .Y(n372) );
  AOI21_X0P7M_A9TR U958 ( .A0(SM14_voltage[5]), .A1(n373), .B0(n372), .Y(n379)
         );
  INV_X0P7M_A9TR U959 ( .A(n374), .Y(n377) );
  AO21A1AI2_X0P7M_A9TR U960 ( .A0(n376), .A1(n379), .B0(n375), .C0(n377), .Y(
        n1069) );
  NOR2B_X1M_A9TR U961 ( .AN(n1069), .B(SM14_voltage[4]), .Y(n378) );
  AOI21_X0P7M_A9TR U962 ( .A0(n380), .A1(SM14_voltage[4]), .B0(n378), .Y(n384)
         );
  NAND2B_X0P5M_A9TR U963 ( .AN(SM14_voltage[3]), .B(n384), .Y(n382) );
  OAI22_X0P5M_A9TR U964 ( .A0(n379), .A1(n378), .B0(SM14_voltage[4]), .B1(n377), .Y(n388) );
  AOI21_X0P7M_A9TR U965 ( .A0(n381), .A1(n1069), .B0(n380), .Y(n386) );
  AOI21_X0P7M_A9TR U966 ( .A0(n382), .A1(n388), .B0(n386), .Y(n1194) );
  XNOR2_X0P7M_A9TR U967 ( .A(SM14_voltage[3]), .B(n1194), .Y(n391) );
  NOR2_X0P7A_A9TR U968 ( .A(SM14_voltage[3]), .B(n1194), .Y(n385) );
  NAND2_X0P5A_A9TR U969 ( .A(n384), .B(n386), .Y(n383) );
  OAI22_X0P5M_A9TR U970 ( .A0(n385), .A1(n384), .B0(n383), .B1(SM14_voltage[3]), .Y(n395) );
  INV_X0P7M_A9TR U971 ( .A(n388), .Y(n387) );
  AOI22_X0P7M_A9TR U972 ( .A0(n388), .A1(n1194), .B0(n387), .B1(n386), .Y(n396) );
  INV_X0P7M_A9TR U973 ( .A(n396), .Y(n389) );
  OA21A1OI2_X0P5M_A9TR U974 ( .A0(SM14_voltage[2]), .A1(n391), .B0(n395), .C0(
        n389), .Y(n393) );
  INV_X0P7M_A9TR U975 ( .A(n393), .Y(n1067) );
  CGENI_X1M_A9TR U976 ( .A(n393), .B(SM14_voltage[1]), .CI(SM14_voltage[2]), 
        .CON(n390) );
  NOR2B_X1M_A9TR U977 ( .AN(n391), .B(n390), .Y(n392) );
  AOI21_X0P7M_A9TR U978 ( .A0(n393), .A1(n395), .B0(n392), .Y(n394) );
  OAI21_X1M_A9TR U979 ( .A0(n396), .A1(n395), .B0(n394), .Y(
        \DUT_controller/N135 ) );
  NOR2_X0P7A_A9TR U980 ( .A(n1067), .B(\DUT_controller/N135 ), .Y(n1195) );
  NOR2_X0P7A_A9TR U981 ( .A(n1194), .B(n1195), .Y(n1193) );
  NOR2_X0P7A_A9TR U982 ( .A(n1193), .B(n1069), .Y(n1068) );
  XNOR2_X0P7M_A9TR U983 ( .A(n1068), .B(n397), .Y(\DUT_controller/N139 ) );
  INV_X0P7M_A9TR U984 ( .A(SM3_voltage[7]), .Y(n399) );
  OAI21_X1M_A9TR U985 ( .A0(n399), .A1(SM3_voltage[5]), .B0(SM3_voltage[6]), 
        .Y(n401) );
  INV_X0P7M_A9TR U986 ( .A(n401), .Y(n407) );
  NOR3_X0P7A_A9TR U987 ( .A(SM3_voltage[5]), .B(SM3_voltage[6]), .C(n399), .Y(
        n400) );
  NOR2_X0P7A_A9TR U988 ( .A(n407), .B(n400), .Y(n406) );
  INV_X0P7M_A9TR U989 ( .A(SM3_voltage[4]), .Y(n402) );
  OAI21_X1M_A9TR U990 ( .A0(SM3_voltage[5]), .A1(SM3_voltage[6]), .B0(
        SM3_voltage[7]), .Y(n423) );
  NOR2_X0P7A_A9TR U991 ( .A(SM3_voltage[5]), .B(n423), .Y(n398) );
  AOI21_X0P7M_A9TR U992 ( .A0(SM3_voltage[5]), .A1(n399), .B0(n398), .Y(n405)
         );
  INV_X0P7M_A9TR U993 ( .A(n400), .Y(n403) );
  AO21A1AI2_X0P7M_A9TR U994 ( .A0(n402), .A1(n405), .B0(n401), .C0(n403), .Y(
        n1097) );
  NOR2B_X1M_A9TR U995 ( .AN(n1097), .B(SM3_voltage[4]), .Y(n404) );
  AOI21_X0P7M_A9TR U996 ( .A0(n406), .A1(SM3_voltage[4]), .B0(n404), .Y(n410)
         );
  NAND2B_X0P5M_A9TR U997 ( .AN(SM3_voltage[3]), .B(n410), .Y(n408) );
  OAI22_X0P5M_A9TR U998 ( .A0(n405), .A1(n404), .B0(SM3_voltage[4]), .B1(n403), 
        .Y(n414) );
  AOI21_X0P7M_A9TR U999 ( .A0(n407), .A1(n1097), .B0(n406), .Y(n412) );
  AOI21_X0P7M_A9TR U1000 ( .A0(n408), .A1(n414), .B0(n412), .Y(n1227) );
  XNOR2_X0P7M_A9TR U1001 ( .A(SM3_voltage[3]), .B(n1227), .Y(n417) );
  NOR2_X0P7A_A9TR U1002 ( .A(SM3_voltage[3]), .B(n1227), .Y(n411) );
  NAND2_X0P5A_A9TR U1003 ( .A(n410), .B(n412), .Y(n409) );
  OAI22_X0P5M_A9TR U1004 ( .A0(n411), .A1(n410), .B0(n409), .B1(SM3_voltage[3]), .Y(n421) );
  INV_X0P7M_A9TR U1005 ( .A(n414), .Y(n413) );
  AOI22_X0P7M_A9TR U1006 ( .A0(n414), .A1(n1227), .B0(n413), .B1(n412), .Y(
        n422) );
  INV_X0P7M_A9TR U1007 ( .A(n422), .Y(n415) );
  OA21A1OI2_X0P5M_A9TR U1008 ( .A0(SM3_voltage[2]), .A1(n417), .B0(n421), .C0(
        n415), .Y(n419) );
  INV_X0P7M_A9TR U1009 ( .A(n419), .Y(n1066) );
  CGENI_X1M_A9TR U1010 ( .A(n419), .B(SM3_voltage[1]), .CI(SM3_voltage[2]), 
        .CON(n416) );
  NOR2B_X1M_A9TR U1011 ( .AN(n417), .B(n416), .Y(n418) );
  AOI21_X0P7M_A9TR U1012 ( .A0(n419), .A1(n421), .B0(n418), .Y(n420) );
  OAI21_X1M_A9TR U1013 ( .A0(n422), .A1(n421), .B0(n420), .Y(
        \DUT_controller/N25 ) );
  NOR2_X0P7A_A9TR U1014 ( .A(n1066), .B(\DUT_controller/N25 ), .Y(n1228) );
  NOR2_X0P7A_A9TR U1015 ( .A(n1227), .B(n1228), .Y(n1226) );
  NOR2_X0P7A_A9TR U1016 ( .A(n1226), .B(n1097), .Y(n1096) );
  XNOR2_X0P7M_A9TR U1017 ( .A(n1096), .B(n423), .Y(\DUT_controller/N29 ) );
  INV_X0P7M_A9TR U1018 ( .A(SM13_voltage[7]), .Y(n425) );
  OAI21_X1M_A9TR U1019 ( .A0(n425), .A1(SM13_voltage[5]), .B0(SM13_voltage[6]), 
        .Y(n427) );
  INV_X0P7M_A9TR U1020 ( .A(n427), .Y(n433) );
  NOR3_X0P7A_A9TR U1021 ( .A(SM13_voltage[5]), .B(SM13_voltage[6]), .C(n425), 
        .Y(n426) );
  NOR2_X0P7A_A9TR U1022 ( .A(n433), .B(n426), .Y(n432) );
  INV_X0P7M_A9TR U1023 ( .A(SM13_voltage[4]), .Y(n428) );
  OAI21_X1M_A9TR U1024 ( .A0(SM13_voltage[5]), .A1(SM13_voltage[6]), .B0(
        SM13_voltage[7]), .Y(n449) );
  NOR2_X0P7A_A9TR U1025 ( .A(SM13_voltage[5]), .B(n449), .Y(n424) );
  AOI21_X0P7M_A9TR U1026 ( .A0(SM13_voltage[5]), .A1(n425), .B0(n424), .Y(n431) );
  INV_X0P7M_A9TR U1027 ( .A(n426), .Y(n429) );
  AO21A1AI2_X0P7M_A9TR U1028 ( .A0(n428), .A1(n431), .B0(n427), .C0(n429), .Y(
        n1074) );
  NOR2B_X1M_A9TR U1029 ( .AN(n1074), .B(SM13_voltage[4]), .Y(n430) );
  AOI21_X0P7M_A9TR U1030 ( .A0(n432), .A1(SM13_voltage[4]), .B0(n430), .Y(n436) );
  NAND2B_X0P5M_A9TR U1031 ( .AN(SM13_voltage[3]), .B(n436), .Y(n434) );
  OAI22_X0P5M_A9TR U1032 ( .A0(n431), .A1(n430), .B0(SM13_voltage[4]), .B1(
        n429), .Y(n440) );
  AOI21_X0P7M_A9TR U1033 ( .A0(n433), .A1(n1074), .B0(n432), .Y(n438) );
  AOI21_X0P7M_A9TR U1034 ( .A0(n434), .A1(n440), .B0(n438), .Y(n1197) );
  XNOR2_X0P7M_A9TR U1035 ( .A(SM13_voltage[3]), .B(n1197), .Y(n443) );
  NOR2_X0P7A_A9TR U1036 ( .A(SM13_voltage[3]), .B(n1197), .Y(n437) );
  NAND2_X0P5A_A9TR U1037 ( .A(n436), .B(n438), .Y(n435) );
  OAI22_X0P5M_A9TR U1038 ( .A0(n437), .A1(n436), .B0(n435), .B1(
        SM13_voltage[3]), .Y(n447) );
  INV_X0P7M_A9TR U1039 ( .A(n440), .Y(n439) );
  AOI22_X0P7M_A9TR U1040 ( .A0(n440), .A1(n1197), .B0(n439), .B1(n438), .Y(
        n448) );
  INV_X0P7M_A9TR U1041 ( .A(n448), .Y(n441) );
  OA21A1OI2_X0P5M_A9TR U1042 ( .A0(SM13_voltage[2]), .A1(n443), .B0(n447), 
        .C0(n441), .Y(n445) );
  INV_X0P7M_A9TR U1043 ( .A(n445), .Y(n1072) );
  CGENI_X1M_A9TR U1044 ( .A(n445), .B(SM13_voltage[1]), .CI(SM13_voltage[2]), 
        .CON(n442) );
  NOR2B_X1M_A9TR U1045 ( .AN(n443), .B(n442), .Y(n444) );
  AOI21_X0P7M_A9TR U1046 ( .A0(n445), .A1(n447), .B0(n444), .Y(n446) );
  OAI21_X1M_A9TR U1047 ( .A0(n448), .A1(n447), .B0(n446), .Y(
        \DUT_controller/N125 ) );
  NOR2_X0P7A_A9TR U1048 ( .A(n1072), .B(\DUT_controller/N125 ), .Y(n1198) );
  NOR2_X0P7A_A9TR U1049 ( .A(n1197), .B(n1198), .Y(n1196) );
  NOR2_X0P7A_A9TR U1050 ( .A(n1196), .B(n1074), .Y(n1073) );
  XNOR2_X0P7M_A9TR U1051 ( .A(n1073), .B(n449), .Y(\DUT_controller/N129 ) );
  INV_X0P7M_A9TR U1052 ( .A(SM4_voltage[7]), .Y(n451) );
  OAI21_X1M_A9TR U1053 ( .A0(n451), .A1(SM4_voltage[5]), .B0(SM4_voltage[6]), 
        .Y(n453) );
  INV_X0P7M_A9TR U1054 ( .A(n453), .Y(n459) );
  NOR3_X0P7A_A9TR U1055 ( .A(SM4_voltage[5]), .B(SM4_voltage[6]), .C(n451), 
        .Y(n452) );
  NOR2_X0P7A_A9TR U1056 ( .A(n459), .B(n452), .Y(n458) );
  INV_X0P7M_A9TR U1057 ( .A(SM4_voltage[4]), .Y(n454) );
  OAI21_X1M_A9TR U1058 ( .A0(SM4_voltage[5]), .A1(SM4_voltage[6]), .B0(
        SM4_voltage[7]), .Y(n475) );
  NOR2_X0P7A_A9TR U1059 ( .A(SM4_voltage[5]), .B(n475), .Y(n450) );
  AOI21_X0P7M_A9TR U1060 ( .A0(SM4_voltage[5]), .A1(n451), .B0(n450), .Y(n457)
         );
  INV_X0P7M_A9TR U1061 ( .A(n452), .Y(n455) );
  AO21A1AI2_X0P7M_A9TR U1062 ( .A0(n454), .A1(n457), .B0(n453), .C0(n455), .Y(
        n1071) );
  NOR2B_X1M_A9TR U1063 ( .AN(n1071), .B(SM4_voltage[4]), .Y(n456) );
  AOI21_X0P7M_A9TR U1064 ( .A0(n458), .A1(SM4_voltage[4]), .B0(n456), .Y(n462)
         );
  NAND2B_X0P5M_A9TR U1065 ( .AN(SM4_voltage[3]), .B(n462), .Y(n460) );
  OAI22_X0P5M_A9TR U1066 ( .A0(n457), .A1(n456), .B0(SM4_voltage[4]), .B1(n455), .Y(n466) );
  AOI21_X0P7M_A9TR U1067 ( .A0(n459), .A1(n1071), .B0(n458), .Y(n464) );
  AOI21_X0P7M_A9TR U1068 ( .A0(n460), .A1(n466), .B0(n464), .Y(n1224) );
  XNOR2_X0P7M_A9TR U1069 ( .A(SM4_voltage[3]), .B(n1224), .Y(n469) );
  NOR2_X0P7A_A9TR U1070 ( .A(SM4_voltage[3]), .B(n1224), .Y(n463) );
  NAND2_X0P5A_A9TR U1071 ( .A(n462), .B(n464), .Y(n461) );
  OAI22_X0P5M_A9TR U1072 ( .A0(n463), .A1(n462), .B0(n461), .B1(SM4_voltage[3]), .Y(n473) );
  INV_X0P7M_A9TR U1073 ( .A(n466), .Y(n465) );
  AOI22_X0P7M_A9TR U1074 ( .A0(n466), .A1(n1224), .B0(n465), .B1(n464), .Y(
        n474) );
  INV_X0P7M_A9TR U1075 ( .A(n474), .Y(n467) );
  OA21A1OI2_X0P5M_A9TR U1076 ( .A0(SM4_voltage[2]), .A1(n469), .B0(n473), .C0(
        n467), .Y(n471) );
  INV_X0P7M_A9TR U1077 ( .A(n471), .Y(n1101) );
  CGENI_X1M_A9TR U1078 ( .A(n471), .B(SM4_voltage[1]), .CI(SM4_voltage[2]), 
        .CON(n468) );
  NOR2B_X1M_A9TR U1079 ( .AN(n469), .B(n468), .Y(n470) );
  AOI21_X0P7M_A9TR U1080 ( .A0(n471), .A1(n473), .B0(n470), .Y(n472) );
  OAI21_X1M_A9TR U1081 ( .A0(n474), .A1(n473), .B0(n472), .Y(
        \DUT_controller/N35 ) );
  NOR2_X0P7A_A9TR U1082 ( .A(n1101), .B(\DUT_controller/N35 ), .Y(n1225) );
  NOR2_X0P7A_A9TR U1083 ( .A(n1224), .B(n1225), .Y(n1223) );
  NOR2_X0P7A_A9TR U1084 ( .A(n1223), .B(n1071), .Y(n1070) );
  XNOR2_X0P7M_A9TR U1085 ( .A(n1070), .B(n475), .Y(\DUT_controller/N39 ) );
  INV_X0P7M_A9TR U1086 ( .A(SM1_voltage[7]), .Y(n477) );
  OAI21_X1M_A9TR U1087 ( .A0(n477), .A1(SM1_voltage[5]), .B0(SM1_voltage[6]), 
        .Y(n479) );
  INV_X0P7M_A9TR U1088 ( .A(n479), .Y(n485) );
  NOR3_X0P7A_A9TR U1089 ( .A(SM1_voltage[5]), .B(SM1_voltage[6]), .C(n477), 
        .Y(n478) );
  NOR2_X0P7A_A9TR U1090 ( .A(n485), .B(n478), .Y(n484) );
  INV_X0P7M_A9TR U1091 ( .A(SM1_voltage[4]), .Y(n480) );
  OAI21_X1M_A9TR U1092 ( .A0(SM1_voltage[5]), .A1(SM1_voltage[6]), .B0(
        SM1_voltage[7]), .Y(n501) );
  NOR2_X0P7A_A9TR U1093 ( .A(SM1_voltage[5]), .B(n501), .Y(n476) );
  AOI21_X0P7M_A9TR U1094 ( .A0(SM1_voltage[5]), .A1(n477), .B0(n476), .Y(n483)
         );
  INV_X0P7M_A9TR U1095 ( .A(n478), .Y(n481) );
  AO21A1AI2_X0P7M_A9TR U1096 ( .A0(n480), .A1(n483), .B0(n479), .C0(n481), .Y(
        n1088) );
  NOR2B_X1M_A9TR U1097 ( .AN(n1088), .B(SM1_voltage[4]), .Y(n482) );
  AOI21_X0P7M_A9TR U1098 ( .A0(n484), .A1(SM1_voltage[4]), .B0(n482), .Y(n488)
         );
  NAND2B_X0P5M_A9TR U1099 ( .AN(SM1_voltage[3]), .B(n488), .Y(n486) );
  OAI22_X0P5M_A9TR U1100 ( .A0(n483), .A1(n482), .B0(SM1_voltage[4]), .B1(n481), .Y(n492) );
  AOI21_X0P7M_A9TR U1101 ( .A0(n485), .A1(n1088), .B0(n484), .Y(n490) );
  AOI21_X0P7M_A9TR U1102 ( .A0(n486), .A1(n492), .B0(n490), .Y(n1233) );
  XNOR2_X0P7M_A9TR U1103 ( .A(SM1_voltage[3]), .B(n1233), .Y(n495) );
  NOR2_X0P7A_A9TR U1104 ( .A(SM1_voltage[3]), .B(n1233), .Y(n489) );
  NAND2_X0P5A_A9TR U1105 ( .A(n488), .B(n490), .Y(n487) );
  OAI22_X0P5M_A9TR U1106 ( .A0(n489), .A1(n488), .B0(n487), .B1(SM1_voltage[3]), .Y(n499) );
  INV_X0P7M_A9TR U1107 ( .A(n492), .Y(n491) );
  AOI22_X0P7M_A9TR U1108 ( .A0(n492), .A1(n1233), .B0(n491), .B1(n490), .Y(
        n500) );
  INV_X0P7M_A9TR U1109 ( .A(n500), .Y(n493) );
  OA21A1OI2_X0P5M_A9TR U1110 ( .A0(SM1_voltage[2]), .A1(n495), .B0(n499), .C0(
        n493), .Y(n497) );
  INV_X0P7M_A9TR U1111 ( .A(n497), .Y(n1086) );
  CGENI_X1M_A9TR U1112 ( .A(n497), .B(SM1_voltage[1]), .CI(SM1_voltage[2]), 
        .CON(n494) );
  NOR2B_X1M_A9TR U1113 ( .AN(n495), .B(n494), .Y(n496) );
  AOI21_X0P7M_A9TR U1114 ( .A0(n497), .A1(n499), .B0(n496), .Y(n498) );
  OAI21_X1M_A9TR U1115 ( .A0(n500), .A1(n499), .B0(n498), .Y(
        \DUT_controller/N5 ) );
  NOR2_X0P7A_A9TR U1116 ( .A(n1086), .B(\DUT_controller/N5 ), .Y(n1234) );
  NOR2_X0P7A_A9TR U1117 ( .A(n1233), .B(n1234), .Y(n1232) );
  NOR2_X0P7A_A9TR U1118 ( .A(n1232), .B(n1088), .Y(n1087) );
  XNOR2_X0P7M_A9TR U1119 ( .A(n1087), .B(n501), .Y(\DUT_controller/N9 ) );
  INV_X0P7M_A9TR U1120 ( .A(SM11_voltage[7]), .Y(n503) );
  OAI21_X1M_A9TR U1121 ( .A0(n503), .A1(SM11_voltage[5]), .B0(SM11_voltage[6]), 
        .Y(n505) );
  INV_X0P7M_A9TR U1122 ( .A(n505), .Y(n511) );
  NOR3_X0P7A_A9TR U1123 ( .A(SM11_voltage[5]), .B(SM11_voltage[6]), .C(n503), 
        .Y(n504) );
  NOR2_X0P7A_A9TR U1124 ( .A(n511), .B(n504), .Y(n510) );
  INV_X0P7M_A9TR U1125 ( .A(SM11_voltage[4]), .Y(n506) );
  OAI21_X1M_A9TR U1126 ( .A0(SM11_voltage[5]), .A1(SM11_voltage[6]), .B0(
        SM11_voltage[7]), .Y(n527) );
  NOR2_X0P7A_A9TR U1127 ( .A(SM11_voltage[5]), .B(n527), .Y(n502) );
  AOI21_X0P7M_A9TR U1128 ( .A0(SM11_voltage[5]), .A1(n503), .B0(n502), .Y(n509) );
  INV_X0P7M_A9TR U1129 ( .A(n504), .Y(n507) );
  AO21A1AI2_X0P7M_A9TR U1130 ( .A0(n506), .A1(n509), .B0(n505), .C0(n507), .Y(
        n1080) );
  NOR2B_X1M_A9TR U1131 ( .AN(n1080), .B(SM11_voltage[4]), .Y(n508) );
  AOI21_X0P7M_A9TR U1132 ( .A0(n510), .A1(SM11_voltage[4]), .B0(n508), .Y(n514) );
  NAND2B_X0P5M_A9TR U1133 ( .AN(SM11_voltage[3]), .B(n514), .Y(n512) );
  OAI22_X0P5M_A9TR U1134 ( .A0(n509), .A1(n508), .B0(SM11_voltage[4]), .B1(
        n507), .Y(n518) );
  AOI21_X0P7M_A9TR U1135 ( .A0(n511), .A1(n1080), .B0(n510), .Y(n516) );
  AOI21_X0P7M_A9TR U1136 ( .A0(n512), .A1(n518), .B0(n516), .Y(n1203) );
  XNOR2_X0P7M_A9TR U1137 ( .A(SM11_voltage[3]), .B(n1203), .Y(n521) );
  NOR2_X0P7A_A9TR U1138 ( .A(SM11_voltage[3]), .B(n1203), .Y(n515) );
  NAND2_X0P5A_A9TR U1139 ( .A(n514), .B(n516), .Y(n513) );
  OAI22_X0P5M_A9TR U1140 ( .A0(n515), .A1(n514), .B0(n513), .B1(
        SM11_voltage[3]), .Y(n525) );
  INV_X0P7M_A9TR U1141 ( .A(n518), .Y(n517) );
  AOI22_X0P7M_A9TR U1142 ( .A0(n518), .A1(n1203), .B0(n517), .B1(n516), .Y(
        n526) );
  INV_X0P7M_A9TR U1143 ( .A(n526), .Y(n519) );
  OA21A1OI2_X0P5M_A9TR U1144 ( .A0(SM11_voltage[2]), .A1(n521), .B0(n525), 
        .C0(n519), .Y(n523) );
  INV_X0P7M_A9TR U1145 ( .A(n523), .Y(n1083) );
  CGENI_X1M_A9TR U1146 ( .A(n523), .B(SM11_voltage[1]), .CI(SM11_voltage[2]), 
        .CON(n520) );
  NOR2B_X1M_A9TR U1147 ( .AN(n521), .B(n520), .Y(n522) );
  AOI21_X0P7M_A9TR U1148 ( .A0(n523), .A1(n525), .B0(n522), .Y(n524) );
  OAI21_X1M_A9TR U1149 ( .A0(n526), .A1(n525), .B0(n524), .Y(
        \DUT_controller/N105 ) );
  NOR2_X0P7A_A9TR U1150 ( .A(n1083), .B(\DUT_controller/N105 ), .Y(n1204) );
  NOR2_X0P7A_A9TR U1151 ( .A(n1203), .B(n1204), .Y(n1202) );
  NOR2_X0P7A_A9TR U1152 ( .A(n1202), .B(n1080), .Y(n1079) );
  XNOR2_X0P7M_A9TR U1153 ( .A(n1079), .B(n527), .Y(\DUT_controller/N109 ) );
  INV_X0P7M_A9TR U1154 ( .A(SM12_voltage[7]), .Y(n529) );
  OAI21_X1M_A9TR U1155 ( .A0(n529), .A1(SM12_voltage[5]), .B0(SM12_voltage[6]), 
        .Y(n531) );
  INV_X0P7M_A9TR U1156 ( .A(n531), .Y(n537) );
  NOR3_X0P7A_A9TR U1157 ( .A(SM12_voltage[5]), .B(SM12_voltage[6]), .C(n529), 
        .Y(n530) );
  NOR2_X0P7A_A9TR U1158 ( .A(n537), .B(n530), .Y(n536) );
  INV_X0P7M_A9TR U1159 ( .A(SM12_voltage[4]), .Y(n532) );
  OAI21_X1M_A9TR U1160 ( .A0(SM12_voltage[5]), .A1(SM12_voltage[6]), .B0(
        SM12_voltage[7]), .Y(n553) );
  NOR2_X0P7A_A9TR U1161 ( .A(SM12_voltage[5]), .B(n553), .Y(n528) );
  AOI21_X0P7M_A9TR U1162 ( .A0(SM12_voltage[5]), .A1(n529), .B0(n528), .Y(n535) );
  INV_X0P7M_A9TR U1163 ( .A(n530), .Y(n533) );
  AO21A1AI2_X0P7M_A9TR U1164 ( .A0(n532), .A1(n535), .B0(n531), .C0(n533), .Y(
        n1082) );
  NOR2B_X1M_A9TR U1165 ( .AN(n1082), .B(SM12_voltage[4]), .Y(n534) );
  AOI21_X0P7M_A9TR U1166 ( .A0(n536), .A1(SM12_voltage[4]), .B0(n534), .Y(n540) );
  NAND2B_X0P5M_A9TR U1167 ( .AN(SM12_voltage[3]), .B(n540), .Y(n538) );
  OAI22_X0P5M_A9TR U1168 ( .A0(n535), .A1(n534), .B0(SM12_voltage[4]), .B1(
        n533), .Y(n544) );
  AOI21_X0P7M_A9TR U1169 ( .A0(n537), .A1(n1082), .B0(n536), .Y(n542) );
  AOI21_X0P7M_A9TR U1170 ( .A0(n538), .A1(n544), .B0(n542), .Y(n1200) );
  XNOR2_X0P7M_A9TR U1171 ( .A(SM12_voltage[3]), .B(n1200), .Y(n547) );
  NOR2_X0P7A_A9TR U1172 ( .A(SM12_voltage[3]), .B(n1200), .Y(n541) );
  NAND2_X0P5A_A9TR U1173 ( .A(n540), .B(n542), .Y(n539) );
  OAI22_X0P5M_A9TR U1174 ( .A0(n541), .A1(n540), .B0(n539), .B1(
        SM12_voltage[3]), .Y(n551) );
  INV_X0P7M_A9TR U1175 ( .A(n544), .Y(n543) );
  AOI22_X0P7M_A9TR U1176 ( .A0(n544), .A1(n1200), .B0(n543), .B1(n542), .Y(
        n552) );
  INV_X0P7M_A9TR U1177 ( .A(n552), .Y(n545) );
  OA21A1OI2_X0P5M_A9TR U1178 ( .A0(SM12_voltage[2]), .A1(n547), .B0(n551), 
        .C0(n545), .Y(n549) );
  INV_X0P7M_A9TR U1179 ( .A(n549), .Y(n1078) );
  CGENI_X1M_A9TR U1180 ( .A(n549), .B(SM12_voltage[1]), .CI(SM12_voltage[2]), 
        .CON(n546) );
  NOR2B_X1M_A9TR U1181 ( .AN(n547), .B(n546), .Y(n548) );
  AOI21_X0P7M_A9TR U1182 ( .A0(n549), .A1(n551), .B0(n548), .Y(n550) );
  OAI21_X1M_A9TR U1183 ( .A0(n552), .A1(n551), .B0(n550), .Y(
        \DUT_controller/N115 ) );
  NOR2_X0P7A_A9TR U1184 ( .A(n1078), .B(\DUT_controller/N115 ), .Y(n1201) );
  NOR2_X0P7A_A9TR U1185 ( .A(n1200), .B(n1201), .Y(n1199) );
  NOR2_X0P7A_A9TR U1186 ( .A(n1199), .B(n1082), .Y(n1081) );
  XNOR2_X0P7M_A9TR U1187 ( .A(n1081), .B(n553), .Y(\DUT_controller/N119 ) );
  INV_X0P7M_A9TR U1188 ( .A(SM9_voltage[7]), .Y(n555) );
  OAI21_X1M_A9TR U1189 ( .A0(n555), .A1(SM9_voltage[5]), .B0(SM9_voltage[6]), 
        .Y(n557) );
  INV_X0P7M_A9TR U1190 ( .A(n557), .Y(n563) );
  NOR3_X0P7A_A9TR U1191 ( .A(SM9_voltage[5]), .B(SM9_voltage[6]), .C(n555), 
        .Y(n556) );
  NOR2_X0P7A_A9TR U1192 ( .A(n563), .B(n556), .Y(n562) );
  INV_X0P7M_A9TR U1193 ( .A(SM9_voltage[4]), .Y(n558) );
  OAI21_X1M_A9TR U1194 ( .A0(SM9_voltage[5]), .A1(SM9_voltage[6]), .B0(
        SM9_voltage[7]), .Y(n579) );
  NOR2_X0P7A_A9TR U1195 ( .A(SM9_voltage[5]), .B(n579), .Y(n554) );
  AOI21_X0P7M_A9TR U1196 ( .A0(SM9_voltage[5]), .A1(n555), .B0(n554), .Y(n561)
         );
  INV_X0P7M_A9TR U1197 ( .A(n556), .Y(n559) );
  AO21A1AI2_X0P7M_A9TR U1198 ( .A0(n558), .A1(n561), .B0(n557), .C0(n559), .Y(
        n1091) );
  NOR2B_X1M_A9TR U1199 ( .AN(n1091), .B(SM9_voltage[4]), .Y(n560) );
  AOI21_X0P7M_A9TR U1200 ( .A0(n562), .A1(SM9_voltage[4]), .B0(n560), .Y(n566)
         );
  NAND2B_X0P5M_A9TR U1201 ( .AN(SM9_voltage[3]), .B(n566), .Y(n564) );
  OAI22_X0P5M_A9TR U1202 ( .A0(n561), .A1(n560), .B0(SM9_voltage[4]), .B1(n559), .Y(n570) );
  AOI21_X0P7M_A9TR U1203 ( .A0(n563), .A1(n1091), .B0(n562), .Y(n568) );
  AOI21_X0P7M_A9TR U1204 ( .A0(n564), .A1(n570), .B0(n568), .Y(n1209) );
  XNOR2_X0P7M_A9TR U1205 ( .A(SM9_voltage[3]), .B(n1209), .Y(n573) );
  NOR2_X0P7A_A9TR U1206 ( .A(SM9_voltage[3]), .B(n1209), .Y(n567) );
  NAND2_X0P5A_A9TR U1207 ( .A(n566), .B(n568), .Y(n565) );
  OAI22_X0P5M_A9TR U1208 ( .A0(n567), .A1(n566), .B0(n565), .B1(SM9_voltage[3]), .Y(n577) );
  INV_X0P7M_A9TR U1209 ( .A(n570), .Y(n569) );
  AOI22_X0P7M_A9TR U1210 ( .A0(n570), .A1(n1209), .B0(n569), .B1(n568), .Y(
        n578) );
  INV_X0P7M_A9TR U1211 ( .A(n578), .Y(n571) );
  OA21A1OI2_X0P5M_A9TR U1212 ( .A0(SM9_voltage[2]), .A1(n573), .B0(n577), .C0(
        n571), .Y(n575) );
  INV_X0P7M_A9TR U1213 ( .A(n575), .Y(n1094) );
  CGENI_X1M_A9TR U1214 ( .A(n575), .B(SM9_voltage[1]), .CI(SM9_voltage[2]), 
        .CON(n572) );
  NOR2B_X1M_A9TR U1215 ( .AN(n573), .B(n572), .Y(n574) );
  AOI21_X0P7M_A9TR U1216 ( .A0(n575), .A1(n577), .B0(n574), .Y(n576) );
  OAI21_X1M_A9TR U1217 ( .A0(n578), .A1(n577), .B0(n576), .Y(
        \DUT_controller/N85 ) );
  NOR2_X0P7A_A9TR U1218 ( .A(n1094), .B(\DUT_controller/N85 ), .Y(n1210) );
  NOR2_X0P7A_A9TR U1219 ( .A(n1209), .B(n1210), .Y(n1208) );
  NOR2_X0P7A_A9TR U1220 ( .A(n1208), .B(n1091), .Y(n1090) );
  XNOR2_X0P7M_A9TR U1221 ( .A(n1090), .B(n579), .Y(\DUT_controller/N89 ) );
  INV_X0P7M_A9TR U1222 ( .A(SM10_voltage[7]), .Y(n581) );
  OAI21_X1M_A9TR U1223 ( .A0(n581), .A1(SM10_voltage[5]), .B0(SM10_voltage[6]), 
        .Y(n583) );
  INV_X0P7M_A9TR U1224 ( .A(n583), .Y(n589) );
  NOR3_X0P7A_A9TR U1225 ( .A(SM10_voltage[5]), .B(SM10_voltage[6]), .C(n581), 
        .Y(n582) );
  NOR2_X0P7A_A9TR U1226 ( .A(n589), .B(n582), .Y(n588) );
  INV_X0P7M_A9TR U1227 ( .A(SM10_voltage[4]), .Y(n584) );
  OAI21_X1M_A9TR U1228 ( .A0(SM10_voltage[5]), .A1(SM10_voltage[6]), .B0(
        SM10_voltage[7]), .Y(n605) );
  NOR2_X0P7A_A9TR U1229 ( .A(SM10_voltage[5]), .B(n605), .Y(n580) );
  AOI21_X0P7M_A9TR U1230 ( .A0(SM10_voltage[5]), .A1(n581), .B0(n580), .Y(n587) );
  INV_X0P7M_A9TR U1231 ( .A(n582), .Y(n585) );
  AO21A1AI2_X0P7M_A9TR U1232 ( .A0(n584), .A1(n587), .B0(n583), .C0(n585), .Y(
        n1085) );
  NOR2B_X1M_A9TR U1233 ( .AN(n1085), .B(SM10_voltage[4]), .Y(n586) );
  AOI21_X0P7M_A9TR U1234 ( .A0(n588), .A1(SM10_voltage[4]), .B0(n586), .Y(n592) );
  NAND2B_X0P5M_A9TR U1235 ( .AN(SM10_voltage[3]), .B(n592), .Y(n590) );
  OAI22_X0P5M_A9TR U1236 ( .A0(n587), .A1(n586), .B0(SM10_voltage[4]), .B1(
        n585), .Y(n596) );
  AOI21_X0P7M_A9TR U1237 ( .A0(n589), .A1(n1085), .B0(n588), .Y(n594) );
  AOI21_X0P7M_A9TR U1238 ( .A0(n590), .A1(n596), .B0(n594), .Y(n1206) );
  XNOR2_X0P7M_A9TR U1239 ( .A(SM10_voltage[3]), .B(n1206), .Y(n599) );
  NOR2_X0P7A_A9TR U1240 ( .A(SM10_voltage[3]), .B(n1206), .Y(n593) );
  NAND2_X0P5A_A9TR U1241 ( .A(n592), .B(n594), .Y(n591) );
  OAI22_X0P5M_A9TR U1242 ( .A0(n593), .A1(n592), .B0(n591), .B1(
        SM10_voltage[3]), .Y(n603) );
  INV_X0P7M_A9TR U1243 ( .A(n596), .Y(n595) );
  AOI22_X0P7M_A9TR U1244 ( .A0(n596), .A1(n1206), .B0(n595), .B1(n594), .Y(
        n604) );
  INV_X0P7M_A9TR U1245 ( .A(n604), .Y(n597) );
  OA21A1OI2_X0P5M_A9TR U1246 ( .A0(SM10_voltage[2]), .A1(n599), .B0(n603), 
        .C0(n597), .Y(n601) );
  INV_X0P7M_A9TR U1247 ( .A(n601), .Y(n1089) );
  CGENI_X1M_A9TR U1248 ( .A(n601), .B(SM10_voltage[1]), .CI(SM10_voltage[2]), 
        .CON(n598) );
  NOR2B_X1M_A9TR U1249 ( .AN(n599), .B(n598), .Y(n600) );
  AOI21_X0P7M_A9TR U1250 ( .A0(n601), .A1(n603), .B0(n600), .Y(n602) );
  OAI21_X1M_A9TR U1251 ( .A0(n604), .A1(n603), .B0(n602), .Y(
        \DUT_controller/N95 ) );
  NOR2_X0P7A_A9TR U1252 ( .A(n1089), .B(\DUT_controller/N95 ), .Y(n1207) );
  NOR2_X0P7A_A9TR U1253 ( .A(n1206), .B(n1207), .Y(n1205) );
  NOR2_X0P7A_A9TR U1254 ( .A(n1205), .B(n1085), .Y(n1084) );
  XNOR2_X0P7M_A9TR U1255 ( .A(n1084), .B(n605), .Y(\DUT_controller/N99 ) );
  INV_X0P7M_A9TR U1256 ( .A(SM2_voltage[7]), .Y(n607) );
  OAI21_X1M_A9TR U1257 ( .A0(n607), .A1(SM2_voltage[5]), .B0(SM2_voltage[6]), 
        .Y(n609) );
  INV_X0P7M_A9TR U1258 ( .A(n609), .Y(n615) );
  NOR3_X0P7A_A9TR U1259 ( .A(SM2_voltage[5]), .B(SM2_voltage[6]), .C(n607), 
        .Y(n608) );
  NOR2_X0P7A_A9TR U1260 ( .A(n615), .B(n608), .Y(n614) );
  INV_X0P7M_A9TR U1261 ( .A(SM2_voltage[4]), .Y(n610) );
  OAI21_X1M_A9TR U1262 ( .A0(SM2_voltage[5]), .A1(SM2_voltage[6]), .B0(
        SM2_voltage[7]), .Y(n631) );
  NOR2_X0P7A_A9TR U1263 ( .A(SM2_voltage[5]), .B(n631), .Y(n606) );
  AOI21_X0P7M_A9TR U1264 ( .A0(SM2_voltage[5]), .A1(n607), .B0(n606), .Y(n613)
         );
  INV_X0P7M_A9TR U1265 ( .A(n608), .Y(n611) );
  AO21A1AI2_X0P7M_A9TR U1266 ( .A0(n610), .A1(n613), .B0(n609), .C0(n611), .Y(
        n1077) );
  NOR2B_X1M_A9TR U1267 ( .AN(n1077), .B(SM2_voltage[4]), .Y(n612) );
  AOI21_X0P7M_A9TR U1268 ( .A0(n614), .A1(SM2_voltage[4]), .B0(n612), .Y(n618)
         );
  NAND2B_X0P5M_A9TR U1269 ( .AN(SM2_voltage[3]), .B(n618), .Y(n616) );
  OAI22_X0P5M_A9TR U1270 ( .A0(n613), .A1(n612), .B0(SM2_voltage[4]), .B1(n611), .Y(n622) );
  AOI21_X0P7M_A9TR U1271 ( .A0(n615), .A1(n1077), .B0(n614), .Y(n620) );
  AOI21_X0P7M_A9TR U1272 ( .A0(n616), .A1(n622), .B0(n620), .Y(n1230) );
  XNOR2_X0P7M_A9TR U1273 ( .A(SM2_voltage[3]), .B(n1230), .Y(n625) );
  NOR2_X0P7A_A9TR U1274 ( .A(SM2_voltage[3]), .B(n1230), .Y(n619) );
  NAND2_X0P5A_A9TR U1275 ( .A(n618), .B(n620), .Y(n617) );
  OAI22_X0P5M_A9TR U1276 ( .A0(n619), .A1(n618), .B0(n617), .B1(SM2_voltage[3]), .Y(n629) );
  INV_X0P7M_A9TR U1277 ( .A(n622), .Y(n621) );
  AOI22_X0P7M_A9TR U1278 ( .A0(n622), .A1(n1230), .B0(n621), .B1(n620), .Y(
        n630) );
  INV_X0P7M_A9TR U1279 ( .A(n630), .Y(n623) );
  OA21A1OI2_X0P5M_A9TR U1280 ( .A0(SM2_voltage[2]), .A1(n625), .B0(n629), .C0(
        n623), .Y(n627) );
  INV_X0P7M_A9TR U1281 ( .A(n627), .Y(n1075) );
  CGENI_X1M_A9TR U1282 ( .A(n627), .B(SM2_voltage[1]), .CI(SM2_voltage[2]), 
        .CON(n624) );
  NOR2B_X1M_A9TR U1283 ( .AN(n625), .B(n624), .Y(n626) );
  AOI21_X0P7M_A9TR U1284 ( .A0(n627), .A1(n629), .B0(n626), .Y(n628) );
  OAI21_X1M_A9TR U1285 ( .A0(n630), .A1(n629), .B0(n628), .Y(
        \DUT_controller/N15 ) );
  NOR2_X0P7A_A9TR U1286 ( .A(n1075), .B(\DUT_controller/N15 ), .Y(n1231) );
  NOR2_X0P7A_A9TR U1287 ( .A(n1230), .B(n1231), .Y(n1229) );
  NOR2_X0P7A_A9TR U1288 ( .A(n1229), .B(n1077), .Y(n1076) );
  XNOR2_X0P7M_A9TR U1289 ( .A(n1076), .B(n631), .Y(\DUT_controller/N19 ) );
  INV_X0P7M_A9TR U1290 ( .A(SM5_voltage[7]), .Y(n633) );
  OAI21_X1M_A9TR U1291 ( .A0(n633), .A1(SM5_voltage[5]), .B0(SM5_voltage[6]), 
        .Y(n635) );
  INV_X0P7M_A9TR U1292 ( .A(n635), .Y(n641) );
  NOR3_X0P7A_A9TR U1293 ( .A(SM5_voltage[5]), .B(SM5_voltage[6]), .C(n633), 
        .Y(n634) );
  NOR2_X0P7A_A9TR U1294 ( .A(n641), .B(n634), .Y(n640) );
  INV_X0P7M_A9TR U1295 ( .A(SM5_voltage[4]), .Y(n636) );
  OAI21_X1M_A9TR U1296 ( .A0(SM5_voltage[5]), .A1(SM5_voltage[6]), .B0(
        SM5_voltage[7]), .Y(n657) );
  NOR2_X0P7A_A9TR U1297 ( .A(SM5_voltage[5]), .B(n657), .Y(n632) );
  AOI21_X0P7M_A9TR U1298 ( .A0(SM5_voltage[5]), .A1(n633), .B0(n632), .Y(n639)
         );
  INV_X0P7M_A9TR U1299 ( .A(n634), .Y(n637) );
  AO21A1AI2_X0P7M_A9TR U1300 ( .A0(n636), .A1(n639), .B0(n635), .C0(n637), .Y(
        n1099) );
  NOR2B_X1M_A9TR U1301 ( .AN(n1099), .B(SM5_voltage[4]), .Y(n638) );
  AOI21_X0P7M_A9TR U1302 ( .A0(n640), .A1(SM5_voltage[4]), .B0(n638), .Y(n644)
         );
  NAND2B_X0P5M_A9TR U1303 ( .AN(SM5_voltage[3]), .B(n644), .Y(n642) );
  OAI22_X0P5M_A9TR U1304 ( .A0(n639), .A1(n638), .B0(SM5_voltage[4]), .B1(n637), .Y(n648) );
  AOI21_X0P7M_A9TR U1305 ( .A0(n641), .A1(n1099), .B0(n640), .Y(n646) );
  AOI21_X0P7M_A9TR U1306 ( .A0(n642), .A1(n648), .B0(n646), .Y(n1221) );
  XNOR2_X0P7M_A9TR U1307 ( .A(SM5_voltage[3]), .B(n1221), .Y(n651) );
  NOR2_X0P7A_A9TR U1308 ( .A(SM5_voltage[3]), .B(n1221), .Y(n645) );
  NAND2_X0P5A_A9TR U1309 ( .A(n644), .B(n646), .Y(n643) );
  OAI22_X0P5M_A9TR U1310 ( .A0(n645), .A1(n644), .B0(n643), .B1(SM5_voltage[3]), .Y(n655) );
  INV_X0P7M_A9TR U1311 ( .A(n648), .Y(n647) );
  AOI22_X0P7M_A9TR U1312 ( .A0(n648), .A1(n1221), .B0(n647), .B1(n646), .Y(
        n656) );
  INV_X0P7M_A9TR U1313 ( .A(n656), .Y(n649) );
  OA21A1OI2_X0P5M_A9TR U1314 ( .A0(SM5_voltage[2]), .A1(n651), .B0(n655), .C0(
        n649), .Y(n653) );
  INV_X0P7M_A9TR U1315 ( .A(n653), .Y(n1100) );
  CGENI_X1M_A9TR U1316 ( .A(n653), .B(SM5_voltage[1]), .CI(SM5_voltage[2]), 
        .CON(n650) );
  NOR2B_X1M_A9TR U1317 ( .AN(n651), .B(n650), .Y(n652) );
  AOI21_X0P7M_A9TR U1318 ( .A0(n653), .A1(n655), .B0(n652), .Y(n654) );
  OAI21_X1M_A9TR U1319 ( .A0(n656), .A1(n655), .B0(n654), .Y(
        \DUT_controller/N45 ) );
  NOR2_X0P7A_A9TR U1320 ( .A(n1100), .B(\DUT_controller/N45 ), .Y(n1222) );
  NOR2_X0P7A_A9TR U1321 ( .A(n1221), .B(n1222), .Y(n1220) );
  NOR2_X0P7A_A9TR U1322 ( .A(n1220), .B(n1099), .Y(n1098) );
  XNOR2_X0P7M_A9TR U1323 ( .A(n1098), .B(n657), .Y(\DUT_controller/N49 ) );
  INV_X0P7M_A9TR U1324 ( .A(SM7_voltage[7]), .Y(n659) );
  OAI21_X1M_A9TR U1325 ( .A0(n659), .A1(SM7_voltage[5]), .B0(SM7_voltage[6]), 
        .Y(n661) );
  INV_X0P7M_A9TR U1326 ( .A(n661), .Y(n667) );
  NOR3_X0P7A_A9TR U1327 ( .A(SM7_voltage[5]), .B(SM7_voltage[6]), .C(n659), 
        .Y(n660) );
  NOR2_X0P7A_A9TR U1328 ( .A(n667), .B(n660), .Y(n666) );
  INV_X0P7M_A9TR U1329 ( .A(SM7_voltage[4]), .Y(n662) );
  OAI21_X1M_A9TR U1330 ( .A0(SM7_voltage[5]), .A1(SM7_voltage[6]), .B0(
        SM7_voltage[7]), .Y(n683) );
  NOR2_X0P7A_A9TR U1331 ( .A(SM7_voltage[5]), .B(n683), .Y(n658) );
  AOI21_X0P7M_A9TR U1332 ( .A0(SM7_voltage[5]), .A1(n659), .B0(n658), .Y(n665)
         );
  INV_X0P7M_A9TR U1333 ( .A(n660), .Y(n663) );
  AO21A1AI2_X0P7M_A9TR U1334 ( .A0(n662), .A1(n665), .B0(n661), .C0(n663), .Y(
        n1059) );
  NOR2B_X1M_A9TR U1335 ( .AN(n1059), .B(SM7_voltage[4]), .Y(n664) );
  AOI21_X0P7M_A9TR U1336 ( .A0(n666), .A1(SM7_voltage[4]), .B0(n664), .Y(n670)
         );
  NAND2B_X0P5M_A9TR U1337 ( .AN(SM7_voltage[3]), .B(n670), .Y(n668) );
  OAI22_X0P5M_A9TR U1338 ( .A0(n665), .A1(n664), .B0(SM7_voltage[4]), .B1(n663), .Y(n674) );
  AOI21_X0P7M_A9TR U1339 ( .A0(n667), .A1(n1059), .B0(n666), .Y(n672) );
  AOI21_X0P7M_A9TR U1340 ( .A0(n668), .A1(n674), .B0(n672), .Y(n1215) );
  XNOR2_X0P7M_A9TR U1341 ( .A(SM7_voltage[3]), .B(n1215), .Y(n677) );
  NOR2_X0P7A_A9TR U1342 ( .A(SM7_voltage[3]), .B(n1215), .Y(n671) );
  NAND2_X0P5A_A9TR U1343 ( .A(n670), .B(n672), .Y(n669) );
  OAI22_X0P5M_A9TR U1344 ( .A0(n671), .A1(n670), .B0(n669), .B1(SM7_voltage[3]), .Y(n681) );
  INV_X0P7M_A9TR U1345 ( .A(n674), .Y(n673) );
  AOI22_X0P7M_A9TR U1346 ( .A0(n674), .A1(n1215), .B0(n673), .B1(n672), .Y(
        n682) );
  INV_X0P7M_A9TR U1347 ( .A(n682), .Y(n675) );
  OA21A1OI2_X0P5M_A9TR U1348 ( .A0(SM7_voltage[2]), .A1(n677), .B0(n681), .C0(
        n675), .Y(n679) );
  INV_X0P7M_A9TR U1349 ( .A(n679), .Y(n1057) );
  CGENI_X1M_A9TR U1350 ( .A(n679), .B(SM7_voltage[1]), .CI(SM7_voltage[2]), 
        .CON(n676) );
  NOR2B_X1M_A9TR U1351 ( .AN(n677), .B(n676), .Y(n678) );
  AOI21_X0P7M_A9TR U1352 ( .A0(n679), .A1(n681), .B0(n678), .Y(n680) );
  OAI21_X1M_A9TR U1353 ( .A0(n682), .A1(n681), .B0(n680), .Y(
        \DUT_controller/N65 ) );
  NOR2_X0P7A_A9TR U1354 ( .A(n1057), .B(\DUT_controller/N65 ), .Y(n1216) );
  NOR2_X0P7A_A9TR U1355 ( .A(n1215), .B(n1216), .Y(n1214) );
  NOR2_X0P7A_A9TR U1356 ( .A(n1214), .B(n1059), .Y(n1058) );
  XNOR2_X0P7M_A9TR U1357 ( .A(n1058), .B(n683), .Y(\DUT_controller/N69 ) );
  INV_X0P7M_A9TR U1358 ( .A(SM6_voltage[7]), .Y(n685) );
  OAI21_X1M_A9TR U1359 ( .A0(n685), .A1(SM6_voltage[5]), .B0(SM6_voltage[6]), 
        .Y(n687) );
  INV_X0P7M_A9TR U1360 ( .A(n687), .Y(n693) );
  NOR3_X0P7A_A9TR U1361 ( .A(SM6_voltage[5]), .B(SM6_voltage[6]), .C(n685), 
        .Y(n686) );
  NOR2_X0P7A_A9TR U1362 ( .A(n693), .B(n686), .Y(n692) );
  INV_X0P7M_A9TR U1363 ( .A(SM6_voltage[4]), .Y(n688) );
  OAI21_X1M_A9TR U1364 ( .A0(SM6_voltage[5]), .A1(SM6_voltage[6]), .B0(
        SM6_voltage[7]), .Y(n709) );
  NOR2_X0P7A_A9TR U1365 ( .A(SM6_voltage[5]), .B(n709), .Y(n684) );
  AOI21_X0P7M_A9TR U1366 ( .A0(SM6_voltage[5]), .A1(n685), .B0(n684), .Y(n691)
         );
  INV_X0P7M_A9TR U1367 ( .A(n686), .Y(n689) );
  AO21A1AI2_X0P7M_A9TR U1368 ( .A0(n688), .A1(n691), .B0(n687), .C0(n689), .Y(
        n1093) );
  NOR2B_X1M_A9TR U1369 ( .AN(n1093), .B(SM6_voltage[4]), .Y(n690) );
  AOI21_X0P7M_A9TR U1370 ( .A0(n692), .A1(SM6_voltage[4]), .B0(n690), .Y(n696)
         );
  NAND2B_X0P5M_A9TR U1371 ( .AN(SM6_voltage[3]), .B(n696), .Y(n694) );
  OAI22_X0P5M_A9TR U1372 ( .A0(n691), .A1(n690), .B0(SM6_voltage[4]), .B1(n689), .Y(n700) );
  AOI21_X0P7M_A9TR U1373 ( .A0(n693), .A1(n1093), .B0(n692), .Y(n698) );
  AOI21_X0P7M_A9TR U1374 ( .A0(n694), .A1(n700), .B0(n698), .Y(n1218) );
  XNOR2_X0P7M_A9TR U1375 ( .A(SM6_voltage[3]), .B(n1218), .Y(n703) );
  NOR2_X0P7A_A9TR U1376 ( .A(SM6_voltage[3]), .B(n1218), .Y(n697) );
  NAND2_X0P5A_A9TR U1377 ( .A(n696), .B(n698), .Y(n695) );
  OAI22_X0P5M_A9TR U1378 ( .A0(n697), .A1(n696), .B0(n695), .B1(SM6_voltage[3]), .Y(n707) );
  INV_X0P7M_A9TR U1379 ( .A(n700), .Y(n699) );
  AOI22_X0P7M_A9TR U1380 ( .A0(n700), .A1(n1218), .B0(n699), .B1(n698), .Y(
        n708) );
  INV_X0P7M_A9TR U1381 ( .A(n708), .Y(n701) );
  OA21A1OI2_X0P5M_A9TR U1382 ( .A0(SM6_voltage[2]), .A1(n703), .B0(n707), .C0(
        n701), .Y(n705) );
  INV_X0P7M_A9TR U1383 ( .A(n705), .Y(n1095) );
  CGENI_X1M_A9TR U1384 ( .A(n705), .B(SM6_voltage[1]), .CI(SM6_voltage[2]), 
        .CON(n702) );
  NOR2B_X1M_A9TR U1385 ( .AN(n703), .B(n702), .Y(n704) );
  AOI21_X0P7M_A9TR U1386 ( .A0(n705), .A1(n707), .B0(n704), .Y(n706) );
  OAI21_X1M_A9TR U1387 ( .A0(n708), .A1(n707), .B0(n706), .Y(
        \DUT_controller/N55 ) );
  NOR2_X0P7A_A9TR U1388 ( .A(n1095), .B(\DUT_controller/N55 ), .Y(n1219) );
  NOR2_X0P7A_A9TR U1389 ( .A(n1218), .B(n1219), .Y(n1217) );
  NOR2_X0P7A_A9TR U1390 ( .A(n1217), .B(n1093), .Y(n1092) );
  XNOR2_X0P7M_A9TR U1391 ( .A(n1092), .B(n709), .Y(\DUT_controller/N59 ) );
  INV_X0P7M_A9TR U1392 ( .A(counter[1]), .Y(n713) );
  NAND2_X0P5A_A9TR U1393 ( .A(n1102), .B(n713), .Y(n712) );
  AND3_X0P7M_A9TR U1394 ( .A(n1102), .B(counter[2]), .C(counter[1]), .Y(n1105)
         );
  NAND2_X0P5A_A9TR U1395 ( .A(n1105), .B(counter[3]), .Y(n1104) );
  XNOR2_X0P7M_A9TR U1396 ( .A(counter[4]), .B(n1104), .Y(N5) );
  NAND2B_X0P5M_A9TR U1397 ( .AN(n1104), .B(counter[4]), .Y(n710) );
  XNOR2_X0P7M_A9TR U1398 ( .A(counter[5]), .B(n710), .Y(N6) );
  NAND4BB_X0P5M_A9TR U1399 ( .AN(counter[2]), .BN(counter[1]), .C(n1102), .D(
        counter[3]), .Y(n711) );
  NOR3_X0P7A_A9TR U1400 ( .A(N5), .B(N6), .C(n711), .Y(n1186) );
  OA21A1OI2_X0P5M_A9TR U1401 ( .A0(n1102), .A1(n713), .B0(n712), .C0(n1186), 
        .Y(N11) );
  NOR2_X0P7A_A9TR U1402 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM1_adjuster/rst [1]), .Y(n1108) );
  AOI211_X0P5M_A9TR U1403 ( .A0(\DUT_SM1_adjuster/rst [1]), .A1(n1102), .B0(
        n1109), .C0(n1108), .Y(n714) );
  INV_X0P7M_A9TR U1404 ( .A(n714), .Y(\DUT_SM1_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1405 ( .A(n1102), .B(\DUT_SM9_adjuster/rst [1]), .Y(n1148)
         );
  AOI211_X0P5M_A9TR U1406 ( .A0(\DUT_SM9_adjuster/rst [1]), .A1(
        \DUT_SM16_adjuster/rst [0]), .B0(n1149), .C0(n1148), .Y(n715) );
  INV_X0P7M_A9TR U1407 ( .A(n715), .Y(\DUT_SM9_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1408 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM10_adjuster/rst [1]), .Y(n1153) );
  AOI211_X0P5M_A9TR U1409 ( .A0(\DUT_SM10_adjuster/rst [1]), .A1(
        \DUT_SM16_adjuster/rst [0]), .B0(n1154), .C0(n1153), .Y(n716) );
  INV_X0P7M_A9TR U1410 ( .A(n716), .Y(\DUT_SM10_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1411 ( .A(n1102), .B(\DUT_SM5_adjuster/rst [1]), .Y(n1128)
         );
  AOI211_X0P5M_A9TR U1412 ( .A0(\DUT_SM5_adjuster/rst [1]), .A1(
        \DUT_SM16_adjuster/rst [0]), .B0(n1129), .C0(n1128), .Y(n717) );
  INV_X0P7M_A9TR U1413 ( .A(n717), .Y(\DUT_SM5_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1414 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM8_adjuster/rst [1]), .Y(n1143) );
  AOI211_X0P5M_A9TR U1415 ( .A0(\DUT_SM8_adjuster/rst [1]), .A1(
        \DUT_SM16_adjuster/rst [0]), .B0(n1144), .C0(n1143), .Y(n718) );
  INV_X0P7M_A9TR U1416 ( .A(n718), .Y(\DUT_SM8_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1417 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM11_adjuster/rst [1]), .Y(n1158) );
  AOI211_X0P5M_A9TR U1418 ( .A0(\DUT_SM11_adjuster/rst [1]), .A1(n1102), .B0(
        n1159), .C0(n1158), .Y(n719) );
  INV_X0P7M_A9TR U1419 ( .A(n719), .Y(\DUT_SM11_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1420 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM12_adjuster/rst [1]), .Y(n1163) );
  AOI211_X0P5M_A9TR U1421 ( .A0(\DUT_SM12_adjuster/rst [1]), .A1(
        \DUT_SM16_adjuster/rst [0]), .B0(n1164), .C0(n1163), .Y(n720) );
  INV_X0P7M_A9TR U1422 ( .A(n720), .Y(\DUT_SM12_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1423 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM13_adjuster/rst [1]), .Y(n1168) );
  AOI211_X0P5M_A9TR U1424 ( .A0(\DUT_SM13_adjuster/rst [1]), .A1(n1102), .B0(
        n1169), .C0(n1168), .Y(n721) );
  INV_X0P7M_A9TR U1425 ( .A(n721), .Y(\DUT_SM13_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1426 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM14_adjuster/rst [1]), .Y(n1173) );
  AOI211_X0P5M_A9TR U1427 ( .A0(\DUT_SM14_adjuster/rst [1]), .A1(
        \DUT_SM16_adjuster/rst [0]), .B0(n1174), .C0(n1173), .Y(n722) );
  INV_X0P7M_A9TR U1428 ( .A(n722), .Y(\DUT_SM14_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1429 ( .A(n1102), .B(\DUT_SM7_adjuster/rst [1]), .Y(n1138)
         );
  AOI211_X0P5M_A9TR U1430 ( .A0(\DUT_SM7_adjuster/rst [1]), .A1(n1102), .B0(
        n1139), .C0(n1138), .Y(n723) );
  INV_X0P7M_A9TR U1431 ( .A(n723), .Y(\DUT_SM7_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1432 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM16_adjuster/rst [1]), .Y(n1182) );
  AOI211_X0P5M_A9TR U1433 ( .A0(\DUT_SM16_adjuster/rst [1]), .A1(n1102), .B0(
        n1183), .C0(n1182), .Y(n724) );
  INV_X0P7M_A9TR U1434 ( .A(n724), .Y(\DUT_SM16_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1435 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM3_adjuster/rst [1]), .Y(n1118) );
  AOI211_X0P5M_A9TR U1436 ( .A0(\DUT_SM3_adjuster/rst [1]), .A1(
        \DUT_SM16_adjuster/rst [0]), .B0(n1119), .C0(n1118), .Y(n725) );
  INV_X0P7M_A9TR U1437 ( .A(n725), .Y(\DUT_SM3_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1438 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM2_adjuster/rst [1]), .Y(n1113) );
  AOI211_X0P5M_A9TR U1439 ( .A0(\DUT_SM2_adjuster/rst [1]), .A1(n1102), .B0(
        n1114), .C0(n1113), .Y(n726) );
  INV_X0P7M_A9TR U1440 ( .A(n726), .Y(\DUT_SM2_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1441 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM4_adjuster/rst [1]), .Y(n1123) );
  AOI211_X0P5M_A9TR U1442 ( .A0(\DUT_SM4_adjuster/rst [1]), .A1(n1102), .B0(
        n1124), .C0(n1123), .Y(n727) );
  INV_X0P7M_A9TR U1443 ( .A(n727), .Y(\DUT_SM4_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1444 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM6_adjuster/rst [1]), .Y(n1133) );
  AOI211_X0P5M_A9TR U1445 ( .A0(\DUT_SM6_adjuster/rst [1]), .A1(
        \DUT_SM16_adjuster/rst [0]), .B0(n1134), .C0(n1133), .Y(n728) );
  INV_X0P7M_A9TR U1446 ( .A(n728), .Y(\DUT_SM6_adjuster/N18 ) );
  NOR2_X0P7A_A9TR U1447 ( .A(\DUT_SM16_adjuster/rst [0]), .B(
        \DUT_SM15_adjuster/rst [1]), .Y(n1178) );
  AOI211_X0P5M_A9TR U1448 ( .A0(\DUT_SM15_adjuster/rst [1]), .A1(
        \DUT_SM16_adjuster/rst [0]), .B0(n1179), .C0(n1178), .Y(n729) );
  INV_X0P7M_A9TR U1449 ( .A(n729), .Y(\DUT_SM15_adjuster/N18 ) );
  AOI22BB_X1M_A9TR U1450 ( .A0(SM7_issued_this_cycle[2]), .A1(n1350), .B0N(
        n1350), .B1N(SM7_issued_this_cycle[2]), .Y(n765) );
  OAI21_X1M_A9TR U1451 ( .A0(n765), .A1(n766), .B0(n1042), .Y(n764) );
  NAND2_X0P5A_A9TR U1452 ( .A(n1139), .B(SM7_issue_width_10_cycle[2]), .Y(n763) );
  AOI22BB_X1M_A9TR U1453 ( .A0(SM8_issued_this_cycle[2]), .A1(n1355), .B0N(
        n1355), .B1N(SM8_issued_this_cycle[2]), .Y(n770) );
  OAI21_X1M_A9TR U1454 ( .A0(n770), .A1(n771), .B0(n1035), .Y(n769) );
  NAND2_X0P5A_A9TR U1455 ( .A(n1144), .B(SM8_issue_width_10_cycle[2]), .Y(n768) );
  AOI22BB_X1M_A9TR U1456 ( .A0(SM9_issued_this_cycle[2]), .A1(n204), .B0N(n204), .B1N(SM9_issued_this_cycle[2]), .Y(n775) );
  OAI21_X1M_A9TR U1457 ( .A0(n775), .A1(n776), .B0(n1028), .Y(n774) );
  NAND2_X0P5A_A9TR U1458 ( .A(n1149), .B(SM9_issue_width_10_cycle[2]), .Y(n773) );
  AOI22BB_X1M_A9TR U1459 ( .A0(SM10_issued_this_cycle[2]), .A1(n1308), .B0N(
        n778), .B1N(SM10_issued_this_cycle[2]), .Y(n781) );
  OAI21_X1M_A9TR U1460 ( .A0(n781), .A1(n782), .B0(n1021), .Y(n780) );
  NAND2_X0P5A_A9TR U1461 ( .A(n1154), .B(SM10_issue_width_10_cycle[2]), .Y(
        n779) );
  AOI22BB_X1M_A9TR U1462 ( .A0(SM11_issued_this_cycle[2]), .A1(n1370), .B0N(
        n1370), .B1N(SM11_issued_this_cycle[2]), .Y(n786) );
  OAI21_X1M_A9TR U1463 ( .A0(n786), .A1(n787), .B0(n1014), .Y(n785) );
  NAND2_X0P5A_A9TR U1464 ( .A(n1159), .B(SM11_issue_width_10_cycle[2]), .Y(
        n784) );
  AOI22BB_X1M_A9TR U1465 ( .A0(SM12_issued_this_cycle[2]), .A1(n1310), .B0N(
        n789), .B1N(SM12_issued_this_cycle[2]), .Y(n792) );
  OAI21_X1M_A9TR U1466 ( .A0(n792), .A1(n793), .B0(n1007), .Y(n791) );
  NAND2_X0P5A_A9TR U1467 ( .A(n1164), .B(SM12_issue_width_10_cycle[2]), .Y(
        n790) );
  AOI22BB_X1M_A9TR U1468 ( .A0(SM13_issued_this_cycle[2]), .A1(n1311), .B0N(
        n795), .B1N(SM13_issued_this_cycle[2]), .Y(n798) );
  OAI21_X1M_A9TR U1469 ( .A0(n798), .A1(n799), .B0(n1000), .Y(n797) );
  NAND2_X0P5A_A9TR U1470 ( .A(n1169), .B(SM13_issue_width_10_cycle[2]), .Y(
        n796) );
  AOI22BB_X1M_A9TR U1471 ( .A0(SM14_issued_this_cycle[2]), .A1(n1385), .B0N(
        n1385), .B1N(SM14_issued_this_cycle[2]), .Y(n803) );
  OAI21_X1M_A9TR U1472 ( .A0(n803), .A1(n804), .B0(n993), .Y(n802) );
  NAND2_X0P5A_A9TR U1473 ( .A(n1174), .B(SM14_issue_width_10_cycle[2]), .Y(
        n801) );
  AOI22BB_X1M_A9TR U1474 ( .A0(SM15_issued_this_cycle[2]), .A1(n1390), .B0N(
        n1390), .B1N(SM15_issued_this_cycle[2]), .Y(n808) );
  OAI21_X1M_A9TR U1475 ( .A0(n808), .A1(n809), .B0(n986), .Y(n807) );
  NAND2_X0P5A_A9TR U1476 ( .A(n1179), .B(SM15_issue_width_10_cycle[2]), .Y(
        n806) );
  AOI22BB_X1M_A9TR U1477 ( .A0(SM16_issued_this_cycle[2]), .A1(n207), .B0N(
        n207), .B1N(SM16_issued_this_cycle[2]), .Y(n813) );
  OAI21_X1M_A9TR U1478 ( .A0(n813), .A1(n814), .B0(n979), .Y(n812) );
  NAND2_X0P5A_A9TR U1479 ( .A(n1183), .B(SM16_issue_width_10_cycle[2]), .Y(
        n811) );
  AOI22BB_X1M_A9TR U1480 ( .A0(SM5_issued_this_cycle[2]), .A1(n202), .B0N(n202), .B1N(SM5_issued_this_cycle[2]), .Y(n818) );
  OAI21_X1M_A9TR U1481 ( .A0(n818), .A1(n819), .B0(n972), .Y(n817) );
  NAND2_X0P5A_A9TR U1482 ( .A(n1129), .B(SM5_issue_width_10_cycle[2]), .Y(n816) );
  AOI22BB_X1M_A9TR U1483 ( .A0(SM6_issued_this_cycle[2]), .A1(n1345), .B0N(
        n1345), .B1N(SM6_issued_this_cycle[2]), .Y(n823) );
  OAI21_X1M_A9TR U1484 ( .A0(n823), .A1(n824), .B0(n965), .Y(n822) );
  NAND2_X0P5A_A9TR U1485 ( .A(n1134), .B(SM6_issue_width_10_cycle[2]), .Y(n821) );
  AOI22BB_X1M_A9TR U1486 ( .A0(SM2_issued_this_cycle[2]), .A1(n1325), .B0N(
        n1325), .B1N(SM2_issued_this_cycle[2]), .Y(n828) );
  OAI21_X1M_A9TR U1487 ( .A0(n828), .A1(n829), .B0(n958), .Y(n827) );
  NAND2_X0P5A_A9TR U1488 ( .A(n1114), .B(SM2_issue_width_10_cycle[2]), .Y(n826) );
  AOI22BB_X1M_A9TR U1489 ( .A0(SM3_issued_this_cycle[2]), .A1(n1330), .B0N(
        n1330), .B1N(SM3_issued_this_cycle[2]), .Y(n833) );
  OAI21_X1M_A9TR U1490 ( .A0(n833), .A1(n834), .B0(n951), .Y(n832) );
  NAND2_X0P5A_A9TR U1491 ( .A(n1119), .B(SM3_issue_width_10_cycle[2]), .Y(n831) );
  AOI22BB_X1M_A9TR U1492 ( .A0(SM4_issued_this_cycle[2]), .A1(n1335), .B0N(
        n1335), .B1N(SM4_issued_this_cycle[2]), .Y(n838) );
  OAI21_X1M_A9TR U1493 ( .A0(n838), .A1(n839), .B0(n944), .Y(n837) );
  NAND2_X0P5A_A9TR U1494 ( .A(n1124), .B(SM4_issue_width_10_cycle[2]), .Y(n836) );
  AOI22BB_X1M_A9TR U1495 ( .A0(SM1_issued_this_cycle[2]), .A1(n1299), .B0N(
        n841), .B1N(SM1_issued_this_cycle[2]), .Y(n844) );
  OAI21_X1M_A9TR U1496 ( .A0(n844), .A1(n845), .B0(n1049), .Y(n843) );
  NAND2_X0P5A_A9TR U1497 ( .A(n1109), .B(SM1_issue_width_10_cycle[2]), .Y(n842) );
  NAND2_X0P5A_A9TR U1498 ( .A(SM13_issued_this_cycle[1]), .B(n847), .Y(n846)
         );
  OAI21_X1M_A9TR U1499 ( .A0(SM13_issued_this_cycle[1]), .A1(n847), .B0(n846), 
        .Y(n850) );
  OAI21_X1M_A9TR U1500 ( .A0(n850), .A1(n851), .B0(n1000), .Y(n849) );
  NAND2_X0P5A_A9TR U1501 ( .A(n1169), .B(SM13_issue_width_10_cycle[1]), .Y(
        n848) );
  NAND2_X0P5A_A9TR U1502 ( .A(SM12_issued_this_cycle[1]), .B(n853), .Y(n852)
         );
  OAI21_X1M_A9TR U1503 ( .A0(SM12_issued_this_cycle[1]), .A1(n853), .B0(n852), 
        .Y(n856) );
  OAI21_X1M_A9TR U1504 ( .A0(n856), .A1(n857), .B0(n1007), .Y(n855) );
  NAND2_X0P5A_A9TR U1505 ( .A(n1164), .B(SM12_issue_width_10_cycle[1]), .Y(
        n854) );
  NAND2_X0P5A_A9TR U1506 ( .A(SM11_issued_this_cycle[1]), .B(n859), .Y(n858)
         );
  OAI21_X1M_A9TR U1507 ( .A0(SM11_issued_this_cycle[1]), .A1(n859), .B0(n858), 
        .Y(n862) );
  OAI21_X1M_A9TR U1508 ( .A0(n862), .A1(n863), .B0(n1014), .Y(n861) );
  NAND2_X0P5A_A9TR U1509 ( .A(n1159), .B(SM11_issue_width_10_cycle[1]), .Y(
        n860) );
  NAND2_X0P5A_A9TR U1510 ( .A(SM10_issued_this_cycle[1]), .B(n865), .Y(n864)
         );
  OAI21_X1M_A9TR U1511 ( .A0(SM10_issued_this_cycle[1]), .A1(n865), .B0(n864), 
        .Y(n868) );
  OAI21_X1M_A9TR U1512 ( .A0(n868), .A1(n869), .B0(n1021), .Y(n867) );
  NAND2_X0P5A_A9TR U1513 ( .A(n1154), .B(SM10_issue_width_10_cycle[1]), .Y(
        n866) );
  NAND2_X0P5A_A9TR U1514 ( .A(SM9_issued_this_cycle[1]), .B(n871), .Y(n870) );
  OAI21_X1M_A9TR U1515 ( .A0(SM9_issued_this_cycle[1]), .A1(n871), .B0(n870), 
        .Y(n874) );
  OAI21_X1M_A9TR U1516 ( .A0(n874), .A1(n875), .B0(n1028), .Y(n873) );
  NAND2_X0P5A_A9TR U1517 ( .A(n1149), .B(SM9_issue_width_10_cycle[1]), .Y(n872) );
  NAND2_X0P5A_A9TR U1518 ( .A(SM8_issued_this_cycle[1]), .B(n877), .Y(n876) );
  OAI21_X1M_A9TR U1519 ( .A0(SM8_issued_this_cycle[1]), .A1(n877), .B0(n876), 
        .Y(n880) );
  OAI21_X1M_A9TR U1520 ( .A0(n880), .A1(n881), .B0(n1035), .Y(n879) );
  NAND2_X0P5A_A9TR U1521 ( .A(n1144), .B(SM8_issue_width_10_cycle[1]), .Y(n878) );
  NAND2_X0P5A_A9TR U1522 ( .A(SM7_issued_this_cycle[1]), .B(n883), .Y(n882) );
  OAI21_X1M_A9TR U1523 ( .A0(SM7_issued_this_cycle[1]), .A1(n883), .B0(n882), 
        .Y(n886) );
  OAI21_X1M_A9TR U1524 ( .A0(n886), .A1(n887), .B0(n1042), .Y(n885) );
  NAND2_X0P5A_A9TR U1525 ( .A(n1139), .B(SM7_issue_width_10_cycle[1]), .Y(n884) );
  NAND2_X0P5A_A9TR U1526 ( .A(SM6_issued_this_cycle[1]), .B(n889), .Y(n888) );
  OAI21_X1M_A9TR U1527 ( .A0(SM6_issued_this_cycle[1]), .A1(n889), .B0(n888), 
        .Y(n892) );
  OAI21_X1M_A9TR U1528 ( .A0(n892), .A1(n893), .B0(n965), .Y(n891) );
  NAND2_X0P5A_A9TR U1529 ( .A(n1134), .B(SM6_issue_width_10_cycle[1]), .Y(n890) );
  NAND2_X0P5A_A9TR U1530 ( .A(SM5_issued_this_cycle[1]), .B(n895), .Y(n894) );
  OAI21_X1M_A9TR U1531 ( .A0(SM5_issued_this_cycle[1]), .A1(n895), .B0(n894), 
        .Y(n898) );
  OAI21_X1M_A9TR U1532 ( .A0(n898), .A1(n899), .B0(n972), .Y(n897) );
  NAND2_X0P5A_A9TR U1533 ( .A(n1129), .B(SM5_issue_width_10_cycle[1]), .Y(n896) );
  NAND2_X0P5A_A9TR U1534 ( .A(SM4_issued_this_cycle[1]), .B(n901), .Y(n900) );
  OAI21_X1M_A9TR U1535 ( .A0(SM4_issued_this_cycle[1]), .A1(n901), .B0(n900), 
        .Y(n904) );
  OAI21_X1M_A9TR U1536 ( .A0(n904), .A1(n905), .B0(n944), .Y(n903) );
  NAND2_X0P5A_A9TR U1537 ( .A(n1124), .B(SM4_issue_width_10_cycle[1]), .Y(n902) );
  NAND2_X0P5A_A9TR U1538 ( .A(SM3_issued_this_cycle[1]), .B(n907), .Y(n906) );
  OAI21_X1M_A9TR U1539 ( .A0(SM3_issued_this_cycle[1]), .A1(n907), .B0(n906), 
        .Y(n910) );
  OAI21_X1M_A9TR U1540 ( .A0(n910), .A1(n911), .B0(n951), .Y(n909) );
  NAND2_X0P5A_A9TR U1541 ( .A(n1119), .B(SM3_issue_width_10_cycle[1]), .Y(n908) );
  NAND2_X0P5A_A9TR U1542 ( .A(SM2_issued_this_cycle[1]), .B(n913), .Y(n912) );
  OAI21_X1M_A9TR U1543 ( .A0(SM2_issued_this_cycle[1]), .A1(n913), .B0(n912), 
        .Y(n916) );
  OAI21_X1M_A9TR U1544 ( .A0(n916), .A1(n917), .B0(n958), .Y(n915) );
  NAND2_X0P5A_A9TR U1545 ( .A(n1114), .B(SM2_issue_width_10_cycle[1]), .Y(n914) );
  NAND2_X0P5A_A9TR U1546 ( .A(SM1_issued_this_cycle[1]), .B(n919), .Y(n918) );
  OAI21_X1M_A9TR U1547 ( .A0(SM1_issued_this_cycle[1]), .A1(n919), .B0(n918), 
        .Y(n922) );
  OAI21_X1M_A9TR U1548 ( .A0(n922), .A1(n923), .B0(n1049), .Y(n921) );
  NAND2_X0P5A_A9TR U1549 ( .A(n1109), .B(SM1_issue_width_10_cycle[1]), .Y(n920) );
  NAND2_X0P5A_A9TR U1550 ( .A(SM15_issued_this_cycle[1]), .B(n925), .Y(n924)
         );
  OAI21_X1M_A9TR U1551 ( .A0(SM15_issued_this_cycle[1]), .A1(n925), .B0(n924), 
        .Y(n928) );
  OAI21_X1M_A9TR U1552 ( .A0(n928), .A1(n929), .B0(n986), .Y(n927) );
  NAND2_X0P5A_A9TR U1553 ( .A(n1179), .B(SM15_issue_width_10_cycle[1]), .Y(
        n926) );
  NAND2_X0P5A_A9TR U1554 ( .A(SM14_issued_this_cycle[1]), .B(n931), .Y(n930)
         );
  OAI21_X1M_A9TR U1555 ( .A0(SM14_issued_this_cycle[1]), .A1(n931), .B0(n930), 
        .Y(n934) );
  OAI21_X1M_A9TR U1556 ( .A0(n934), .A1(n935), .B0(n993), .Y(n933) );
  NAND2_X0P5A_A9TR U1557 ( .A(n1174), .B(SM14_issue_width_10_cycle[1]), .Y(
        n932) );
  NAND2_X0P5A_A9TR U1558 ( .A(SM16_issued_this_cycle[1]), .B(n937), .Y(n936)
         );
  OAI21_X1M_A9TR U1559 ( .A0(SM16_issued_this_cycle[1]), .A1(n937), .B0(n936), 
        .Y(n940) );
  OAI21_X1M_A9TR U1560 ( .A0(n940), .A1(n941), .B0(n979), .Y(n939) );
  NAND2_X0P5A_A9TR U1561 ( .A(n1183), .B(SM16_issue_width_10_cycle[1]), .Y(
        n938) );
  NAND2_X0P5A_A9TR U1562 ( .A(SM4_issued_this_cycle[3]), .B(n943), .Y(n942) );
  OAI21_X1M_A9TR U1563 ( .A0(SM4_issued_this_cycle[3]), .A1(n943), .B0(n942), 
        .Y(n947) );
  OAI21_X1M_A9TR U1564 ( .A0(n947), .A1(n948), .B0(n944), .Y(n946) );
  NAND2_X0P5A_A9TR U1565 ( .A(n1124), .B(SM4_issue_width_10_cycle[3]), .Y(n945) );
  NAND2_X0P5A_A9TR U1566 ( .A(SM3_issued_this_cycle[3]), .B(n950), .Y(n949) );
  OAI21_X1M_A9TR U1567 ( .A0(SM3_issued_this_cycle[3]), .A1(n950), .B0(n949), 
        .Y(n954) );
  OAI21_X1M_A9TR U1568 ( .A0(n954), .A1(n955), .B0(n951), .Y(n953) );
  NAND2_X0P5A_A9TR U1569 ( .A(n1119), .B(SM3_issue_width_10_cycle[3]), .Y(n952) );
  NAND2_X0P5A_A9TR U1570 ( .A(SM2_issued_this_cycle[3]), .B(n957), .Y(n956) );
  OAI21_X1M_A9TR U1571 ( .A0(SM2_issued_this_cycle[3]), .A1(n957), .B0(n956), 
        .Y(n961) );
  OAI21_X1M_A9TR U1572 ( .A0(n961), .A1(n962), .B0(n958), .Y(n960) );
  NAND2_X0P5A_A9TR U1573 ( .A(n1114), .B(SM2_issue_width_10_cycle[3]), .Y(n959) );
  NAND2_X0P5A_A9TR U1574 ( .A(SM6_issued_this_cycle[3]), .B(n964), .Y(n963) );
  OAI21_X1M_A9TR U1575 ( .A0(SM6_issued_this_cycle[3]), .A1(n964), .B0(n963), 
        .Y(n968) );
  OAI21_X1M_A9TR U1576 ( .A0(n968), .A1(n969), .B0(n965), .Y(n967) );
  NAND2_X0P5A_A9TR U1577 ( .A(n1134), .B(SM6_issue_width_10_cycle[3]), .Y(n966) );
  NAND2_X0P5A_A9TR U1578 ( .A(SM5_issued_this_cycle[3]), .B(n971), .Y(n970) );
  OAI21_X1M_A9TR U1579 ( .A0(SM5_issued_this_cycle[3]), .A1(n971), .B0(n970), 
        .Y(n975) );
  OAI21_X1M_A9TR U1580 ( .A0(n975), .A1(n976), .B0(n972), .Y(n974) );
  NAND2_X0P5A_A9TR U1581 ( .A(n1129), .B(SM5_issue_width_10_cycle[3]), .Y(n973) );
  NAND2_X0P5A_A9TR U1582 ( .A(SM16_issued_this_cycle[3]), .B(n978), .Y(n977)
         );
  OAI21_X1M_A9TR U1583 ( .A0(SM16_issued_this_cycle[3]), .A1(n978), .B0(n977), 
        .Y(n982) );
  OAI21_X1M_A9TR U1584 ( .A0(n982), .A1(n983), .B0(n979), .Y(n981) );
  NAND2_X0P5A_A9TR U1585 ( .A(n1183), .B(SM16_issue_width_10_cycle[3]), .Y(
        n980) );
  NAND2_X0P5A_A9TR U1586 ( .A(SM15_issued_this_cycle[3]), .B(n985), .Y(n984)
         );
  OAI21_X1M_A9TR U1587 ( .A0(SM15_issued_this_cycle[3]), .A1(n985), .B0(n984), 
        .Y(n989) );
  OAI21_X1M_A9TR U1588 ( .A0(n989), .A1(n990), .B0(n986), .Y(n988) );
  NAND2_X0P5A_A9TR U1589 ( .A(n1179), .B(SM15_issue_width_10_cycle[3]), .Y(
        n987) );
  NAND2_X0P5A_A9TR U1590 ( .A(SM14_issued_this_cycle[3]), .B(n992), .Y(n991)
         );
  OAI21_X1M_A9TR U1591 ( .A0(SM14_issued_this_cycle[3]), .A1(n992), .B0(n991), 
        .Y(n996) );
  OAI21_X1M_A9TR U1592 ( .A0(n996), .A1(n997), .B0(n993), .Y(n995) );
  NAND2_X0P5A_A9TR U1593 ( .A(n1174), .B(SM14_issue_width_10_cycle[3]), .Y(
        n994) );
  NAND2_X0P5A_A9TR U1594 ( .A(SM13_issued_this_cycle[3]), .B(n999), .Y(n998)
         );
  OAI21_X1M_A9TR U1595 ( .A0(SM13_issued_this_cycle[3]), .A1(n999), .B0(n998), 
        .Y(n1003) );
  OAI21_X1M_A9TR U1596 ( .A0(n1003), .A1(n1004), .B0(n1000), .Y(n1002) );
  NAND2_X0P5A_A9TR U1597 ( .A(n1169), .B(SM13_issue_width_10_cycle[3]), .Y(
        n1001) );
  NAND2_X0P5A_A9TR U1598 ( .A(SM12_issued_this_cycle[3]), .B(n1006), .Y(n1005)
         );
  OAI21_X1M_A9TR U1599 ( .A0(SM12_issued_this_cycle[3]), .A1(n1006), .B0(n1005), .Y(n1010) );
  OAI21_X1M_A9TR U1600 ( .A0(n1010), .A1(n1011), .B0(n1007), .Y(n1009) );
  NAND2_X0P5A_A9TR U1601 ( .A(n1164), .B(SM12_issue_width_10_cycle[3]), .Y(
        n1008) );
  NAND2_X0P5A_A9TR U1602 ( .A(SM11_issued_this_cycle[3]), .B(n1013), .Y(n1012)
         );
  OAI21_X1M_A9TR U1603 ( .A0(SM11_issued_this_cycle[3]), .A1(n1013), .B0(n1012), .Y(n1017) );
  OAI21_X1M_A9TR U1604 ( .A0(n1017), .A1(n1018), .B0(n1014), .Y(n1016) );
  NAND2_X0P5A_A9TR U1605 ( .A(n1159), .B(SM11_issue_width_10_cycle[3]), .Y(
        n1015) );
  NAND2_X0P5A_A9TR U1606 ( .A(SM10_issued_this_cycle[3]), .B(n1020), .Y(n1019)
         );
  OAI21_X1M_A9TR U1607 ( .A0(SM10_issued_this_cycle[3]), .A1(n1020), .B0(n1019), .Y(n1024) );
  OAI21_X1M_A9TR U1608 ( .A0(n1024), .A1(n1025), .B0(n1021), .Y(n1023) );
  NAND2_X0P5A_A9TR U1609 ( .A(n1154), .B(SM10_issue_width_10_cycle[3]), .Y(
        n1022) );
  NAND2_X0P5A_A9TR U1610 ( .A(SM9_issued_this_cycle[3]), .B(n1027), .Y(n1026)
         );
  OAI21_X1M_A9TR U1611 ( .A0(SM9_issued_this_cycle[3]), .A1(n1027), .B0(n1026), 
        .Y(n1031) );
  OAI21_X1M_A9TR U1612 ( .A0(n1031), .A1(n1032), .B0(n1028), .Y(n1030) );
  NAND2_X0P5A_A9TR U1613 ( .A(n1149), .B(SM9_issue_width_10_cycle[3]), .Y(
        n1029) );
  NAND2_X0P5A_A9TR U1614 ( .A(SM8_issued_this_cycle[3]), .B(n1034), .Y(n1033)
         );
  OAI21_X1M_A9TR U1615 ( .A0(SM8_issued_this_cycle[3]), .A1(n1034), .B0(n1033), 
        .Y(n1038) );
  OAI21_X1M_A9TR U1616 ( .A0(n1038), .A1(n1039), .B0(n1035), .Y(n1037) );
  NAND2_X0P5A_A9TR U1617 ( .A(n1144), .B(SM8_issue_width_10_cycle[3]), .Y(
        n1036) );
  NAND2_X0P5A_A9TR U1618 ( .A(SM7_issued_this_cycle[3]), .B(n1041), .Y(n1040)
         );
  OAI21_X1M_A9TR U1619 ( .A0(SM7_issued_this_cycle[3]), .A1(n1041), .B0(n1040), 
        .Y(n1045) );
  OAI21_X1M_A9TR U1620 ( .A0(n1045), .A1(n1046), .B0(n1042), .Y(n1044) );
  NAND2_X0P5A_A9TR U1621 ( .A(n1139), .B(SM7_issue_width_10_cycle[3]), .Y(
        n1043) );
  NAND2_X0P5A_A9TR U1622 ( .A(SM1_issued_this_cycle[3]), .B(n1048), .Y(n1047)
         );
  OAI21_X1M_A9TR U1623 ( .A0(SM1_issued_this_cycle[3]), .A1(n1048), .B0(n1047), 
        .Y(n1052) );
  OAI21_X1M_A9TR U1624 ( .A0(n1052), .A1(n1053), .B0(n1049), .Y(n1051) );
  NAND2_X0P5A_A9TR U1625 ( .A(n1109), .B(SM1_issue_width_10_cycle[3]), .Y(
        n1050) );
  AOI21_X0P7M_A9TR U1626 ( .A0(n1054), .A1(\DUT_controller/N75 ), .B0(n1213), 
        .Y(\DUT_controller/N76 ) );
  AOI21_X0P7M_A9TR U1627 ( .A0(n1211), .A1(n1056), .B0(n1055), .Y(
        \DUT_controller/N78 ) );
  AOI21_X0P7M_A9TR U1628 ( .A0(n1057), .A1(\DUT_controller/N65 ), .B0(n1216), 
        .Y(\DUT_controller/N66 ) );
  AOI21_X0P7M_A9TR U1629 ( .A0(n1214), .A1(n1059), .B0(n1058), .Y(
        \DUT_controller/N68 ) );
  AOI21_X0P7M_A9TR U1630 ( .A0(n1060), .A1(\DUT_controller/N155 ), .B0(n1189), 
        .Y(\DUT_controller/N156 ) );
  AOI21_X0P7M_A9TR U1631 ( .A0(n1187), .A1(n1062), .B0(n1061), .Y(
        \DUT_controller/N158 ) );
  AOI21_X0P7M_A9TR U1632 ( .A0(n1063), .A1(\DUT_controller/N145 ), .B0(n1192), 
        .Y(\DUT_controller/N146 ) );
  AOI21_X0P7M_A9TR U1633 ( .A0(n1190), .A1(n1065), .B0(n1064), .Y(
        \DUT_controller/N148 ) );
  AOI21_X0P7M_A9TR U1634 ( .A0(n1066), .A1(\DUT_controller/N25 ), .B0(n1228), 
        .Y(\DUT_controller/N26 ) );
  AOI21_X0P7M_A9TR U1635 ( .A0(n1067), .A1(\DUT_controller/N135 ), .B0(n1195), 
        .Y(\DUT_controller/N136 ) );
  AOI21_X0P7M_A9TR U1636 ( .A0(n1193), .A1(n1069), .B0(n1068), .Y(
        \DUT_controller/N138 ) );
  AOI21_X0P7M_A9TR U1637 ( .A0(n1223), .A1(n1071), .B0(n1070), .Y(
        \DUT_controller/N38 ) );
  AOI21_X0P7M_A9TR U1638 ( .A0(n1072), .A1(\DUT_controller/N125 ), .B0(n1198), 
        .Y(\DUT_controller/N126 ) );
  AOI21_X0P7M_A9TR U1639 ( .A0(n1196), .A1(n1074), .B0(n1073), .Y(
        \DUT_controller/N128 ) );
  AOI21_X0P7M_A9TR U1640 ( .A0(n1075), .A1(\DUT_controller/N15 ), .B0(n1231), 
        .Y(\DUT_controller/N16 ) );
  AOI21_X0P7M_A9TR U1641 ( .A0(n1229), .A1(n1077), .B0(n1076), .Y(
        \DUT_controller/N18 ) );
  AOI21_X0P7M_A9TR U1642 ( .A0(n1078), .A1(\DUT_controller/N115 ), .B0(n1201), 
        .Y(\DUT_controller/N116 ) );
  AOI21_X0P7M_A9TR U1643 ( .A0(n1202), .A1(n1080), .B0(n1079), .Y(
        \DUT_controller/N108 ) );
  AOI21_X0P7M_A9TR U1644 ( .A0(n1199), .A1(n1082), .B0(n1081), .Y(
        \DUT_controller/N118 ) );
  AOI21_X0P7M_A9TR U1645 ( .A0(n1083), .A1(\DUT_controller/N105 ), .B0(n1204), 
        .Y(\DUT_controller/N106 ) );
  AOI21_X0P7M_A9TR U1646 ( .A0(n1205), .A1(n1085), .B0(n1084), .Y(
        \DUT_controller/N98 ) );
  AOI21_X0P7M_A9TR U1647 ( .A0(n1086), .A1(\DUT_controller/N5 ), .B0(n1234), 
        .Y(\DUT_controller/N6 ) );
  AOI21_X0P7M_A9TR U1648 ( .A0(n1232), .A1(n1088), .B0(n1087), .Y(
        \DUT_controller/N8 ) );
  AOI21_X0P7M_A9TR U1649 ( .A0(n1089), .A1(\DUT_controller/N95 ), .B0(n1207), 
        .Y(\DUT_controller/N96 ) );
  AOI21_X0P7M_A9TR U1650 ( .A0(n1208), .A1(n1091), .B0(n1090), .Y(
        \DUT_controller/N88 ) );
  AOI21_X0P7M_A9TR U1651 ( .A0(n1217), .A1(n1093), .B0(n1092), .Y(
        \DUT_controller/N58 ) );
  AOI21_X0P7M_A9TR U1652 ( .A0(n1094), .A1(\DUT_controller/N85 ), .B0(n1210), 
        .Y(\DUT_controller/N86 ) );
  AOI21_X0P7M_A9TR U1653 ( .A0(n1095), .A1(\DUT_controller/N55 ), .B0(n1219), 
        .Y(\DUT_controller/N56 ) );
  AOI21_X0P7M_A9TR U1654 ( .A0(n1226), .A1(n1097), .B0(n1096), .Y(
        \DUT_controller/N28 ) );
  AOI21_X0P7M_A9TR U1655 ( .A0(n1220), .A1(n1099), .B0(n1098), .Y(
        \DUT_controller/N48 ) );
  AOI21_X0P7M_A9TR U1656 ( .A0(n1100), .A1(\DUT_controller/N45 ), .B0(n1222), 
        .Y(\DUT_controller/N46 ) );
  AOI21_X0P7M_A9TR U1657 ( .A0(n1101), .A1(\DUT_controller/N35 ), .B0(n1225), 
        .Y(\DUT_controller/N36 ) );
  AOI21_X0P7M_A9TR U1658 ( .A0(n1102), .A1(counter[1]), .B0(counter[2]), .Y(
        n1103) );
  NOR2_X0P7A_A9TR U1659 ( .A(n1105), .B(n1103), .Y(N3) );
  OAI21_X1M_A9TR U1660 ( .A0(n1105), .A1(counter[3]), .B0(n1104), .Y(n1106) );
  NOR2_X0P7A_A9TR U1661 ( .A(n1186), .B(n1106), .Y(N13) );
  NAND2_X0P5A_A9TR U1662 ( .A(n1108), .B(n1107), .Y(n1111) );
  OAI21_X1M_A9TR U1663 ( .A0(n1108), .A1(n1107), .B0(n1111), .Y(
        \DUT_SM1_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1664 ( .A0(\DUT_SM1_adjuster/rst [3]), .A1(n1111), .B0(
        n1109), .Y(n1110) );
  OAI21_X1M_A9TR U1665 ( .A0(\DUT_SM1_adjuster/rst [3]), .A1(n1111), .B0(n1110), .Y(\DUT_SM1_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1666 ( .A(n1113), .B(n1112), .Y(n1116) );
  OAI21_X1M_A9TR U1667 ( .A0(n1113), .A1(n1112), .B0(n1116), .Y(
        \DUT_SM2_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1668 ( .A0(\DUT_SM2_adjuster/rst [3]), .A1(n1116), .B0(
        n1114), .Y(n1115) );
  OAI21_X1M_A9TR U1669 ( .A0(\DUT_SM2_adjuster/rst [3]), .A1(n1116), .B0(n1115), .Y(\DUT_SM2_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1670 ( .A(n1118), .B(n1117), .Y(n1121) );
  OAI21_X1M_A9TR U1671 ( .A0(n1118), .A1(n1117), .B0(n1121), .Y(
        \DUT_SM3_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1672 ( .A0(\DUT_SM3_adjuster/rst [3]), .A1(n1121), .B0(
        n1119), .Y(n1120) );
  OAI21_X1M_A9TR U1673 ( .A0(\DUT_SM3_adjuster/rst [3]), .A1(n1121), .B0(n1120), .Y(\DUT_SM3_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1674 ( .A(n1123), .B(n1122), .Y(n1126) );
  OAI21_X1M_A9TR U1675 ( .A0(n1123), .A1(n1122), .B0(n1126), .Y(
        \DUT_SM4_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1676 ( .A0(\DUT_SM4_adjuster/rst [3]), .A1(n1126), .B0(
        n1124), .Y(n1125) );
  OAI21_X1M_A9TR U1677 ( .A0(\DUT_SM4_adjuster/rst [3]), .A1(n1126), .B0(n1125), .Y(\DUT_SM4_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1678 ( .A(n1128), .B(n1127), .Y(n1131) );
  OAI21_X1M_A9TR U1679 ( .A0(n1128), .A1(n1127), .B0(n1131), .Y(
        \DUT_SM5_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1680 ( .A0(\DUT_SM5_adjuster/rst [3]), .A1(n1131), .B0(
        n1129), .Y(n1130) );
  OAI21_X1M_A9TR U1681 ( .A0(\DUT_SM5_adjuster/rst [3]), .A1(n1131), .B0(n1130), .Y(\DUT_SM5_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1682 ( .A(n1133), .B(n1132), .Y(n1136) );
  OAI21_X1M_A9TR U1683 ( .A0(n1133), .A1(n1132), .B0(n1136), .Y(
        \DUT_SM6_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1684 ( .A0(\DUT_SM6_adjuster/rst [3]), .A1(n1136), .B0(
        n1134), .Y(n1135) );
  OAI21_X1M_A9TR U1685 ( .A0(\DUT_SM6_adjuster/rst [3]), .A1(n1136), .B0(n1135), .Y(\DUT_SM6_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1686 ( .A(n1138), .B(n1137), .Y(n1141) );
  OAI21_X1M_A9TR U1687 ( .A0(n1138), .A1(n1137), .B0(n1141), .Y(
        \DUT_SM7_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1688 ( .A0(\DUT_SM7_adjuster/rst [3]), .A1(n1141), .B0(
        n1139), .Y(n1140) );
  OAI21_X1M_A9TR U1689 ( .A0(\DUT_SM7_adjuster/rst [3]), .A1(n1141), .B0(n1140), .Y(\DUT_SM7_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1690 ( .A(n1143), .B(n1142), .Y(n1146) );
  OAI21_X1M_A9TR U1691 ( .A0(n1143), .A1(n1142), .B0(n1146), .Y(
        \DUT_SM8_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1692 ( .A0(\DUT_SM8_adjuster/rst [3]), .A1(n1146), .B0(
        n1144), .Y(n1145) );
  OAI21_X1M_A9TR U1693 ( .A0(\DUT_SM8_adjuster/rst [3]), .A1(n1146), .B0(n1145), .Y(\DUT_SM8_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1694 ( .A(n1148), .B(n1147), .Y(n1151) );
  OAI21_X1M_A9TR U1695 ( .A0(n1148), .A1(n1147), .B0(n1151), .Y(
        \DUT_SM9_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1696 ( .A0(\DUT_SM9_adjuster/rst [3]), .A1(n1151), .B0(
        n1149), .Y(n1150) );
  OAI21_X1M_A9TR U1697 ( .A0(\DUT_SM9_adjuster/rst [3]), .A1(n1151), .B0(n1150), .Y(\DUT_SM9_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1698 ( .A(n1153), .B(n1152), .Y(n1156) );
  OAI21_X1M_A9TR U1699 ( .A0(n1153), .A1(n1152), .B0(n1156), .Y(
        \DUT_SM10_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1700 ( .A0(\DUT_SM10_adjuster/rst [3]), .A1(n1156), .B0(
        n1154), .Y(n1155) );
  OAI21_X1M_A9TR U1701 ( .A0(\DUT_SM10_adjuster/rst [3]), .A1(n1156), .B0(
        n1155), .Y(\DUT_SM10_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1702 ( .A(n1158), .B(n1157), .Y(n1161) );
  OAI21_X1M_A9TR U1703 ( .A0(n1158), .A1(n1157), .B0(n1161), .Y(
        \DUT_SM11_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1704 ( .A0(\DUT_SM11_adjuster/rst [3]), .A1(n1161), .B0(
        n1159), .Y(n1160) );
  OAI21_X1M_A9TR U1705 ( .A0(\DUT_SM11_adjuster/rst [3]), .A1(n1161), .B0(
        n1160), .Y(\DUT_SM11_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1706 ( .A(n1163), .B(n1162), .Y(n1166) );
  OAI21_X1M_A9TR U1707 ( .A0(n1163), .A1(n1162), .B0(n1166), .Y(
        \DUT_SM12_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1708 ( .A0(\DUT_SM12_adjuster/rst [3]), .A1(n1166), .B0(
        n1164), .Y(n1165) );
  OAI21_X1M_A9TR U1709 ( .A0(\DUT_SM12_adjuster/rst [3]), .A1(n1166), .B0(
        n1165), .Y(\DUT_SM12_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1710 ( .A(n1168), .B(n1167), .Y(n1171) );
  OAI21_X1M_A9TR U1711 ( .A0(n1168), .A1(n1167), .B0(n1171), .Y(
        \DUT_SM13_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1712 ( .A0(\DUT_SM13_adjuster/rst [3]), .A1(n1171), .B0(
        n1169), .Y(n1170) );
  OAI21_X1M_A9TR U1713 ( .A0(\DUT_SM13_adjuster/rst [3]), .A1(n1171), .B0(
        n1170), .Y(\DUT_SM13_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1714 ( .A(n1173), .B(n1172), .Y(n1176) );
  OAI21_X1M_A9TR U1715 ( .A0(n1173), .A1(n1172), .B0(n1176), .Y(
        \DUT_SM14_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1716 ( .A0(\DUT_SM14_adjuster/rst [3]), .A1(n1176), .B0(
        n1174), .Y(n1175) );
  OAI21_X1M_A9TR U1717 ( .A0(\DUT_SM14_adjuster/rst [3]), .A1(n1176), .B0(
        n1175), .Y(\DUT_SM14_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1718 ( .A(n1178), .B(n1177), .Y(n1181) );
  OAI21_X1M_A9TR U1719 ( .A0(n1178), .A1(n1177), .B0(n1181), .Y(
        \DUT_SM15_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1720 ( .A0(\DUT_SM15_adjuster/rst [3]), .A1(n1181), .B0(
        n1179), .Y(n1180) );
  OAI21_X1M_A9TR U1721 ( .A0(\DUT_SM15_adjuster/rst [3]), .A1(n1181), .B0(
        n1180), .Y(\DUT_SM15_adjuster/N20 ) );
  NAND2_X0P5A_A9TR U1722 ( .A(n1182), .B(n1316), .Y(n1185) );
  OAI21_X1M_A9TR U1723 ( .A0(n1182), .A1(n1316), .B0(n1185), .Y(
        \DUT_SM16_adjuster/N19 ) );
  AOI21_X0P7M_A9TR U1724 ( .A0(\DUT_SM16_adjuster/rst [3]), .A1(n1185), .B0(
        n1183), .Y(n1184) );
  OAI21_X1M_A9TR U1725 ( .A0(\DUT_SM16_adjuster/rst [3]), .A1(n1185), .B0(
        n1184), .Y(\DUT_SM16_adjuster/N20 ) );
  XOR2_X0P7M_A9TR U1726 ( .A(clk_controller), .B(n1186), .Y(n195) );
  AO21_X1M_A9TR U1727 ( .A0(n1189), .A1(n1188), .B0(n1187), .Y(
        \DUT_controller/N157 ) );
  AO21_X1M_A9TR U1728 ( .A0(n1192), .A1(n1191), .B0(n1190), .Y(
        \DUT_controller/N147 ) );
  AO21_X1M_A9TR U1729 ( .A0(n1195), .A1(n1194), .B0(n1193), .Y(
        \DUT_controller/N137 ) );
  AO21_X1M_A9TR U1730 ( .A0(n1198), .A1(n1197), .B0(n1196), .Y(
        \DUT_controller/N127 ) );
  AO21_X1M_A9TR U1731 ( .A0(n1201), .A1(n1200), .B0(n1199), .Y(
        \DUT_controller/N117 ) );
  AO21_X1M_A9TR U1732 ( .A0(n1204), .A1(n1203), .B0(n1202), .Y(
        \DUT_controller/N107 ) );
  AO21_X1M_A9TR U1733 ( .A0(n1207), .A1(n1206), .B0(n1205), .Y(
        \DUT_controller/N97 ) );
  AO21_X1M_A9TR U1734 ( .A0(n1210), .A1(n1209), .B0(n1208), .Y(
        \DUT_controller/N87 ) );
  AO21_X1M_A9TR U1735 ( .A0(n1213), .A1(n1212), .B0(n1211), .Y(
        \DUT_controller/N77 ) );
  AO21_X1M_A9TR U1736 ( .A0(n1216), .A1(n1215), .B0(n1214), .Y(
        \DUT_controller/N67 ) );
  AO21_X1M_A9TR U1737 ( .A0(n1219), .A1(n1218), .B0(n1217), .Y(
        \DUT_controller/N57 ) );
  AO21_X1M_A9TR U1738 ( .A0(n1222), .A1(n1221), .B0(n1220), .Y(
        \DUT_controller/N47 ) );
  AO21_X1M_A9TR U1739 ( .A0(n1225), .A1(n1224), .B0(n1223), .Y(
        \DUT_controller/N37 ) );
  AO21_X1M_A9TR U1740 ( .A0(n1228), .A1(n1227), .B0(n1226), .Y(
        \DUT_controller/N27 ) );
  AO21_X1M_A9TR U1741 ( .A0(n1231), .A1(n1230), .B0(n1229), .Y(
        \DUT_controller/N17 ) );
  AO21_X1M_A9TR U1742 ( .A0(n1234), .A1(n1233), .B0(n1232), .Y(
        \DUT_controller/N7 ) );
endmodule

